module TLMonitor_54( // @[:freechips.rocketchip.system.DefaultConfig.fir@219780.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultConfig.fir@219781.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultConfig.fir@219782.4]
  input         io_in_a_ready, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input         io_in_a_valid, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [2:0]  io_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [2:0]  io_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [2:0]  io_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [5:0]  io_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [32:0] io_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [7:0]  io_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input         io_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input         io_in_d_ready, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input         io_in_d_valid, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [2:0]  io_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [2:0]  io_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
  input  [5:0]  io_in_d_bits_source // @[:freechips.rocketchip.system.DefaultConfig.fir@219783.4]
);
  wire [31:0] plusarg_reader_out; // @[PlusArg.scala 42:11:freechips.rocketchip.system.DefaultConfig.fir@220930.4]
  wire [12:0] _T_36; // @[package.scala 185:77:freechips.rocketchip.system.DefaultConfig.fir@219810.6]
  wire [5:0] _T_37; // @[package.scala 185:82:freechips.rocketchip.system.DefaultConfig.fir@219811.6]
  wire [5:0] _T_38; // @[package.scala 185:46:freechips.rocketchip.system.DefaultConfig.fir@219812.6]
  wire [32:0] _GEN_18; // @[Edges.scala 21:16:freechips.rocketchip.system.DefaultConfig.fir@219813.6]
  wire [32:0] _T_39; // @[Edges.scala 21:16:freechips.rocketchip.system.DefaultConfig.fir@219813.6]
  wire  _T_40; // @[Edges.scala 21:24:freechips.rocketchip.system.DefaultConfig.fir@219814.6]
  wire [1:0] _T_42; // @[OneHot.scala 51:49:freechips.rocketchip.system.DefaultConfig.fir@219816.6]
  wire [3:0] _T_43; // @[OneHot.scala 52:12:freechips.rocketchip.system.DefaultConfig.fir@219817.6]
  wire [2:0] _T_44; // @[OneHot.scala 52:27:freechips.rocketchip.system.DefaultConfig.fir@219818.6]
  wire [2:0] _T_45; // @[Misc.scala 206:81:freechips.rocketchip.system.DefaultConfig.fir@219819.6]
  wire  _T_46; // @[Misc.scala 210:21:freechips.rocketchip.system.DefaultConfig.fir@219820.6]
  wire  _T_47; // @[Misc.scala 213:26:freechips.rocketchip.system.DefaultConfig.fir@219821.6]
  wire  _T_48; // @[Misc.scala 214:26:freechips.rocketchip.system.DefaultConfig.fir@219822.6]
  wire  _T_49; // @[Misc.scala 215:20:freechips.rocketchip.system.DefaultConfig.fir@219823.6]
  wire  _T_51; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219825.6]
  wire  _T_52; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219826.6]
  wire  _T_54; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219828.6]
  wire  _T_55; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219829.6]
  wire  _T_56; // @[Misc.scala 213:26:freechips.rocketchip.system.DefaultConfig.fir@219830.6]
  wire  _T_57; // @[Misc.scala 214:26:freechips.rocketchip.system.DefaultConfig.fir@219831.6]
  wire  _T_58; // @[Misc.scala 215:20:freechips.rocketchip.system.DefaultConfig.fir@219832.6]
  wire  _T_59; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219833.6]
  wire  _T_60; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219834.6]
  wire  _T_61; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219835.6]
  wire  _T_62; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219836.6]
  wire  _T_63; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219837.6]
  wire  _T_64; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219838.6]
  wire  _T_65; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219839.6]
  wire  _T_66; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219840.6]
  wire  _T_67; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219841.6]
  wire  _T_68; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219842.6]
  wire  _T_69; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219843.6]
  wire  _T_70; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219844.6]
  wire  _T_71; // @[Misc.scala 213:26:freechips.rocketchip.system.DefaultConfig.fir@219845.6]
  wire  _T_72; // @[Misc.scala 214:26:freechips.rocketchip.system.DefaultConfig.fir@219846.6]
  wire  _T_73; // @[Misc.scala 215:20:freechips.rocketchip.system.DefaultConfig.fir@219847.6]
  wire  _T_74; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219848.6]
  wire  _T_75; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219849.6]
  wire  _T_76; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219850.6]
  wire  _T_77; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219851.6]
  wire  _T_78; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219852.6]
  wire  _T_79; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219853.6]
  wire  _T_80; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219854.6]
  wire  _T_81; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219855.6]
  wire  _T_82; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219856.6]
  wire  _T_83; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219857.6]
  wire  _T_84; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219858.6]
  wire  _T_85; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219859.6]
  wire  _T_86; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219860.6]
  wire  _T_87; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219861.6]
  wire  _T_88; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219862.6]
  wire  _T_89; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219863.6]
  wire  _T_90; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219864.6]
  wire  _T_91; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219865.6]
  wire  _T_92; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219866.6]
  wire  _T_93; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219867.6]
  wire  _T_94; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219868.6]
  wire  _T_95; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219869.6]
  wire  _T_96; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219870.6]
  wire  _T_97; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219871.6]
  wire [1:0] _T_98; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219872.6]
  wire [1:0] _T_99; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219873.6]
  wire [3:0] _T_100; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219874.6]
  wire [1:0] _T_101; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219875.6]
  wire [1:0] _T_102; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219876.6]
  wire [3:0] _T_103; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219877.6]
  wire [7:0] _T_104; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219878.6]
  wire  _T_105; // @[Monitor.scala 40:25:freechips.rocketchip.system.DefaultConfig.fir@219879.6]
  wire [32:0] _T_107; // @[Parameters.scala 121:31:freechips.rocketchip.system.DefaultConfig.fir@219882.8]
  wire [33:0] _T_108; // @[Parameters.scala 121:49:freechips.rocketchip.system.DefaultConfig.fir@219883.8]
  wire [33:0] _T_109; // @[Parameters.scala 121:52:freechips.rocketchip.system.DefaultConfig.fir@219884.8]
  wire [33:0] _T_110; // @[Parameters.scala 121:52:freechips.rocketchip.system.DefaultConfig.fir@219885.8]
  wire  _T_111; // @[Parameters.scala 121:67:freechips.rocketchip.system.DefaultConfig.fir@219886.8]
  wire  _T_116; // @[Monitor.scala 41:14:freechips.rocketchip.system.DefaultConfig.fir@219891.8]
  wire  _T_125; // @[Monitor.scala 44:14:freechips.rocketchip.system.DefaultConfig.fir@219912.8]
  wire  _T_126; // @[Monitor.scala 44:14:freechips.rocketchip.system.DefaultConfig.fir@219913.8]
  wire  _T_128; // @[Monitor.scala 45:14:freechips.rocketchip.system.DefaultConfig.fir@219919.8]
  wire  _T_129; // @[Monitor.scala 45:14:freechips.rocketchip.system.DefaultConfig.fir@219920.8]
  wire  _T_130; // @[Bundles.scala 109:27:freechips.rocketchip.system.DefaultConfig.fir@219925.8]
  wire  _T_132; // @[Monitor.scala 46:14:freechips.rocketchip.system.DefaultConfig.fir@219927.8]
  wire  _T_133; // @[Monitor.scala 46:14:freechips.rocketchip.system.DefaultConfig.fir@219928.8]
  wire [7:0] _T_134; // @[Monitor.scala 47:15:freechips.rocketchip.system.DefaultConfig.fir@219933.8]
  wire  _T_135; // @[Monitor.scala 47:28:freechips.rocketchip.system.DefaultConfig.fir@219934.8]
  wire  _T_137; // @[Monitor.scala 47:14:freechips.rocketchip.system.DefaultConfig.fir@219936.8]
  wire  _T_138; // @[Monitor.scala 47:14:freechips.rocketchip.system.DefaultConfig.fir@219937.8]
  wire  _T_139; // @[Monitor.scala 48:15:freechips.rocketchip.system.DefaultConfig.fir@219942.8]
  wire  _T_141; // @[Monitor.scala 48:14:freechips.rocketchip.system.DefaultConfig.fir@219944.8]
  wire  _T_142; // @[Monitor.scala 48:14:freechips.rocketchip.system.DefaultConfig.fir@219945.8]
  wire  _T_143; // @[Monitor.scala 51:25:freechips.rocketchip.system.DefaultConfig.fir@219951.6]
  wire  _T_172; // @[Monitor.scala 58:28:freechips.rocketchip.system.DefaultConfig.fir@220005.8]
  wire  _T_174; // @[Monitor.scala 58:14:freechips.rocketchip.system.DefaultConfig.fir@220007.8]
  wire  _T_175; // @[Monitor.scala 58:14:freechips.rocketchip.system.DefaultConfig.fir@220008.8]
  wire  _T_185; // @[Monitor.scala 63:25:freechips.rocketchip.system.DefaultConfig.fir@220031.6]
  wire  _T_187; // @[Parameters.scala 90:42:freechips.rocketchip.system.DefaultConfig.fir@220034.8]
  wire  _T_195; // @[Parameters.scala 168:56:freechips.rocketchip.system.DefaultConfig.fir@220042.8]
  wire  _T_198; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220045.8]
  wire  _T_199; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220046.8]
  wire  _T_206; // @[Monitor.scala 67:28:freechips.rocketchip.system.DefaultConfig.fir@220065.8]
  wire  _T_208; // @[Monitor.scala 67:14:freechips.rocketchip.system.DefaultConfig.fir@220067.8]
  wire  _T_209; // @[Monitor.scala 67:14:freechips.rocketchip.system.DefaultConfig.fir@220068.8]
  wire  _T_210; // @[Monitor.scala 68:27:freechips.rocketchip.system.DefaultConfig.fir@220073.8]
  wire  _T_212; // @[Monitor.scala 68:14:freechips.rocketchip.system.DefaultConfig.fir@220075.8]
  wire  _T_213; // @[Monitor.scala 68:14:freechips.rocketchip.system.DefaultConfig.fir@220076.8]
  wire  _T_218; // @[Monitor.scala 72:25:freechips.rocketchip.system.DefaultConfig.fir@220090.6]
  wire  _T_247; // @[Monitor.scala 80:25:freechips.rocketchip.system.DefaultConfig.fir@220141.6]
  wire [7:0] _T_272; // @[Monitor.scala 85:30:freechips.rocketchip.system.DefaultConfig.fir@220183.8]
  wire [7:0] _T_273; // @[Monitor.scala 85:28:freechips.rocketchip.system.DefaultConfig.fir@220184.8]
  wire  _T_274; // @[Monitor.scala 85:37:freechips.rocketchip.system.DefaultConfig.fir@220185.8]
  wire  _T_276; // @[Monitor.scala 85:14:freechips.rocketchip.system.DefaultConfig.fir@220187.8]
  wire  _T_277; // @[Monitor.scala 85:14:freechips.rocketchip.system.DefaultConfig.fir@220188.8]
  wire  _T_278; // @[Monitor.scala 88:25:freechips.rocketchip.system.DefaultConfig.fir@220194.6]
  wire  _T_296; // @[Bundles.scala 139:33:freechips.rocketchip.system.DefaultConfig.fir@220225.8]
  wire  _T_298; // @[Monitor.scala 92:14:freechips.rocketchip.system.DefaultConfig.fir@220227.8]
  wire  _T_299; // @[Monitor.scala 92:14:freechips.rocketchip.system.DefaultConfig.fir@220228.8]
  wire  _T_304; // @[Monitor.scala 96:25:freechips.rocketchip.system.DefaultConfig.fir@220242.6]
  wire  _T_322; // @[Bundles.scala 146:30:freechips.rocketchip.system.DefaultConfig.fir@220273.8]
  wire  _T_324; // @[Monitor.scala 100:14:freechips.rocketchip.system.DefaultConfig.fir@220275.8]
  wire  _T_325; // @[Monitor.scala 100:14:freechips.rocketchip.system.DefaultConfig.fir@220276.8]
  wire  _T_330; // @[Monitor.scala 104:25:freechips.rocketchip.system.DefaultConfig.fir@220290.6]
  wire  _T_356; // @[Bundles.scala 43:24:freechips.rocketchip.system.DefaultConfig.fir@220340.6]
  wire  _T_358; // @[Monitor.scala 256:12:freechips.rocketchip.system.DefaultConfig.fir@220342.6]
  wire  _T_359; // @[Monitor.scala 256:12:freechips.rocketchip.system.DefaultConfig.fir@220343.6]
  wire  _T_376; // @[Monitor.scala 263:25:freechips.rocketchip.system.DefaultConfig.fir@220360.6]
  wire  _T_380; // @[Monitor.scala 265:27:freechips.rocketchip.system.DefaultConfig.fir@220369.8]
  wire  _T_382; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220371.8]
  wire  _T_383; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220372.8]
  wire  _T_396; // @[Monitor.scala 271:25:freechips.rocketchip.system.DefaultConfig.fir@220402.6]
  wire  _T_424; // @[Monitor.scala 281:25:freechips.rocketchip.system.DefaultConfig.fir@220460.6]
  wire  _T_517; // @[Bundles.scala 283:22:freechips.rocketchip.system.DefaultConfig.fir@220650.4]
  wire [2:0] _T_522; // @[Edges.scala 220:59:freechips.rocketchip.system.DefaultConfig.fir@220655.4]
  wire  _T_523; // @[Edges.scala 92:37:freechips.rocketchip.system.DefaultConfig.fir@220656.4]
  wire  _T_524; // @[Edges.scala 92:28:freechips.rocketchip.system.DefaultConfig.fir@220657.4]
  reg [2:0] _T_527; // @[Edges.scala 229:27:freechips.rocketchip.system.DefaultConfig.fir@220659.4]
  reg [31:0] _RAND_0;
  wire [3:0] _T_528; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220660.4]
  wire [3:0] _T_529; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220661.4]
  wire [2:0] _T_530; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220662.4]
  wire  _T_531; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220663.4]
  reg [2:0] _T_540; // @[Monitor.scala 337:22:freechips.rocketchip.system.DefaultConfig.fir@220674.4]
  reg [31:0] _RAND_1;
  reg [2:0] _T_542; // @[Monitor.scala 338:22:freechips.rocketchip.system.DefaultConfig.fir@220675.4]
  reg [31:0] _RAND_2;
  reg [2:0] _T_544; // @[Monitor.scala 339:22:freechips.rocketchip.system.DefaultConfig.fir@220676.4]
  reg [31:0] _RAND_3;
  reg [5:0] _T_546; // @[Monitor.scala 340:22:freechips.rocketchip.system.DefaultConfig.fir@220677.4]
  reg [31:0] _RAND_4;
  reg [32:0] _T_548; // @[Monitor.scala 341:22:freechips.rocketchip.system.DefaultConfig.fir@220678.4]
  reg [63:0] _RAND_5;
  wire  _T_549; // @[Monitor.scala 342:22:freechips.rocketchip.system.DefaultConfig.fir@220679.4]
  wire  _T_550; // @[Monitor.scala 342:19:freechips.rocketchip.system.DefaultConfig.fir@220680.4]
  wire  _T_551; // @[Monitor.scala 343:29:freechips.rocketchip.system.DefaultConfig.fir@220682.6]
  wire  _T_553; // @[Monitor.scala 343:14:freechips.rocketchip.system.DefaultConfig.fir@220684.6]
  wire  _T_554; // @[Monitor.scala 343:14:freechips.rocketchip.system.DefaultConfig.fir@220685.6]
  wire  _T_555; // @[Monitor.scala 344:29:freechips.rocketchip.system.DefaultConfig.fir@220690.6]
  wire  _T_557; // @[Monitor.scala 344:14:freechips.rocketchip.system.DefaultConfig.fir@220692.6]
  wire  _T_558; // @[Monitor.scala 344:14:freechips.rocketchip.system.DefaultConfig.fir@220693.6]
  wire  _T_559; // @[Monitor.scala 345:29:freechips.rocketchip.system.DefaultConfig.fir@220698.6]
  wire  _T_561; // @[Monitor.scala 345:14:freechips.rocketchip.system.DefaultConfig.fir@220700.6]
  wire  _T_562; // @[Monitor.scala 345:14:freechips.rocketchip.system.DefaultConfig.fir@220701.6]
  wire  _T_563; // @[Monitor.scala 346:29:freechips.rocketchip.system.DefaultConfig.fir@220706.6]
  wire  _T_565; // @[Monitor.scala 346:14:freechips.rocketchip.system.DefaultConfig.fir@220708.6]
  wire  _T_566; // @[Monitor.scala 346:14:freechips.rocketchip.system.DefaultConfig.fir@220709.6]
  wire  _T_567; // @[Monitor.scala 347:29:freechips.rocketchip.system.DefaultConfig.fir@220714.6]
  wire  _T_569; // @[Monitor.scala 347:14:freechips.rocketchip.system.DefaultConfig.fir@220716.6]
  wire  _T_570; // @[Monitor.scala 347:14:freechips.rocketchip.system.DefaultConfig.fir@220717.6]
  wire  _T_572; // @[Monitor.scala 349:20:freechips.rocketchip.system.DefaultConfig.fir@220724.4]
  wire  _T_573; // @[Bundles.scala 283:22:freechips.rocketchip.system.DefaultConfig.fir@220732.4]
  wire [12:0] _T_575; // @[package.scala 185:77:freechips.rocketchip.system.DefaultConfig.fir@220734.4]
  wire [5:0] _T_576; // @[package.scala 185:82:freechips.rocketchip.system.DefaultConfig.fir@220735.4]
  wire [5:0] _T_577; // @[package.scala 185:46:freechips.rocketchip.system.DefaultConfig.fir@220736.4]
  wire [2:0] _T_578; // @[Edges.scala 220:59:freechips.rocketchip.system.DefaultConfig.fir@220737.4]
  wire  _T_579; // @[Edges.scala 106:36:freechips.rocketchip.system.DefaultConfig.fir@220738.4]
  reg [2:0] _T_582; // @[Edges.scala 229:27:freechips.rocketchip.system.DefaultConfig.fir@220740.4]
  reg [31:0] _RAND_6;
  wire [3:0] _T_583; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220741.4]
  wire [3:0] _T_584; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220742.4]
  wire [2:0] _T_585; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220743.4]
  wire  _T_586; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220744.4]
  reg [2:0] _T_595; // @[Monitor.scala 406:22:freechips.rocketchip.system.DefaultConfig.fir@220755.4]
  reg [31:0] _RAND_7;
  reg [2:0] _T_599; // @[Monitor.scala 408:22:freechips.rocketchip.system.DefaultConfig.fir@220757.4]
  reg [31:0] _RAND_8;
  reg [5:0] _T_601; // @[Monitor.scala 409:22:freechips.rocketchip.system.DefaultConfig.fir@220758.4]
  reg [31:0] _RAND_9;
  wire  _T_606; // @[Monitor.scala 412:22:freechips.rocketchip.system.DefaultConfig.fir@220761.4]
  wire  _T_607; // @[Monitor.scala 412:19:freechips.rocketchip.system.DefaultConfig.fir@220762.4]
  wire  _T_608; // @[Monitor.scala 413:29:freechips.rocketchip.system.DefaultConfig.fir@220764.6]
  wire  _T_610; // @[Monitor.scala 413:14:freechips.rocketchip.system.DefaultConfig.fir@220766.6]
  wire  _T_611; // @[Monitor.scala 413:14:freechips.rocketchip.system.DefaultConfig.fir@220767.6]
  wire  _T_616; // @[Monitor.scala 415:29:freechips.rocketchip.system.DefaultConfig.fir@220780.6]
  wire  _T_618; // @[Monitor.scala 415:14:freechips.rocketchip.system.DefaultConfig.fir@220782.6]
  wire  _T_619; // @[Monitor.scala 415:14:freechips.rocketchip.system.DefaultConfig.fir@220783.6]
  wire  _T_620; // @[Monitor.scala 416:29:freechips.rocketchip.system.DefaultConfig.fir@220788.6]
  wire  _T_622; // @[Monitor.scala 416:14:freechips.rocketchip.system.DefaultConfig.fir@220790.6]
  wire  _T_623; // @[Monitor.scala 416:14:freechips.rocketchip.system.DefaultConfig.fir@220791.6]
  wire  _T_633; // @[Monitor.scala 420:20:freechips.rocketchip.system.DefaultConfig.fir@220814.4]
  reg [63:0] _T_635; // @[Monitor.scala 440:27:freechips.rocketchip.system.DefaultConfig.fir@220823.4]
  reg [63:0] _RAND_10;
  reg [2:0] _T_646; // @[Edges.scala 229:27:freechips.rocketchip.system.DefaultConfig.fir@220833.4]
  reg [31:0] _RAND_11;
  wire [3:0] _T_647; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220834.4]
  wire [3:0] _T_648; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220835.4]
  wire [2:0] _T_649; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220836.4]
  wire  _T_650; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220837.4]
  reg [2:0] _T_667; // @[Edges.scala 229:27:freechips.rocketchip.system.DefaultConfig.fir@220856.4]
  reg [31:0] _RAND_12;
  wire [3:0] _T_668; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220857.4]
  wire [3:0] _T_669; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220858.4]
  wire [2:0] _T_670; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220859.4]
  wire  _T_671; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220860.4]
  wire  _T_682; // @[Monitor.scala 446:27:freechips.rocketchip.system.DefaultConfig.fir@220875.4]
  wire [63:0] _T_684; // @[OneHot.scala 45:35:freechips.rocketchip.system.DefaultConfig.fir@220878.6]
  wire [63:0] _T_685; // @[Monitor.scala 448:23:freechips.rocketchip.system.DefaultConfig.fir@220880.6]
  wire  _T_686; // @[Monitor.scala 448:23:freechips.rocketchip.system.DefaultConfig.fir@220881.6]
  wire  _T_687; // @[Monitor.scala 448:14:freechips.rocketchip.system.DefaultConfig.fir@220882.6]
  wire  _T_689; // @[Monitor.scala 448:13:freechips.rocketchip.system.DefaultConfig.fir@220884.6]
  wire  _T_690; // @[Monitor.scala 448:13:freechips.rocketchip.system.DefaultConfig.fir@220885.6]
  wire [63:0] _GEN_15; // @[Monitor.scala 446:72:freechips.rocketchip.system.DefaultConfig.fir@220877.4]
  wire  _T_695; // @[Monitor.scala 453:27:freechips.rocketchip.system.DefaultConfig.fir@220896.4]
  wire  _T_697; // @[Monitor.scala 453:75:freechips.rocketchip.system.DefaultConfig.fir@220898.4]
  wire  _T_698; // @[Monitor.scala 453:72:freechips.rocketchip.system.DefaultConfig.fir@220899.4]
  wire [63:0] _T_699; // @[OneHot.scala 45:35:freechips.rocketchip.system.DefaultConfig.fir@220901.6]
  wire [63:0] _T_700; // @[Monitor.scala 455:21:freechips.rocketchip.system.DefaultConfig.fir@220903.6]
  wire [63:0] _T_701; // @[Monitor.scala 455:32:freechips.rocketchip.system.DefaultConfig.fir@220904.6]
  wire  _T_702; // @[Monitor.scala 455:32:freechips.rocketchip.system.DefaultConfig.fir@220905.6]
  wire  _T_704; // @[Monitor.scala 455:13:freechips.rocketchip.system.DefaultConfig.fir@220907.6]
  wire  _T_705; // @[Monitor.scala 455:13:freechips.rocketchip.system.DefaultConfig.fir@220908.6]
  wire [63:0] _GEN_16; // @[Monitor.scala 453:91:freechips.rocketchip.system.DefaultConfig.fir@220900.4]
  wire  _T_706; // @[Monitor.scala 459:20:freechips.rocketchip.system.DefaultConfig.fir@220914.4]
  wire  _T_707; // @[Monitor.scala 459:40:freechips.rocketchip.system.DefaultConfig.fir@220915.4]
  wire  _T_708; // @[Monitor.scala 459:33:freechips.rocketchip.system.DefaultConfig.fir@220916.4]
  wire  _T_709; // @[Monitor.scala 459:30:freechips.rocketchip.system.DefaultConfig.fir@220917.4]
  wire  _T_711; // @[Monitor.scala 459:13:freechips.rocketchip.system.DefaultConfig.fir@220919.4]
  wire  _T_712; // @[Monitor.scala 459:13:freechips.rocketchip.system.DefaultConfig.fir@220920.4]
  wire [63:0] _T_713; // @[Monitor.scala 462:27:freechips.rocketchip.system.DefaultConfig.fir@220925.4]
  wire [63:0] _T_714; // @[Monitor.scala 462:38:freechips.rocketchip.system.DefaultConfig.fir@220926.4]
  wire [63:0] _T_715; // @[Monitor.scala 462:36:freechips.rocketchip.system.DefaultConfig.fir@220927.4]
  reg [31:0] _T_717; // @[Monitor.scala 464:27:freechips.rocketchip.system.DefaultConfig.fir@220929.4]
  reg [31:0] _RAND_13;
  wire  _T_718; // @[Monitor.scala 467:23:freechips.rocketchip.system.DefaultConfig.fir@220932.4]
  wire  _T_719; // @[Monitor.scala 467:13:freechips.rocketchip.system.DefaultConfig.fir@220933.4]
  wire  _T_720; // @[Monitor.scala 467:36:freechips.rocketchip.system.DefaultConfig.fir@220934.4]
  wire  _T_721; // @[Monitor.scala 467:27:freechips.rocketchip.system.DefaultConfig.fir@220935.4]
  wire  _T_722; // @[Monitor.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@220936.4]
  wire  _T_723; // @[Monitor.scala 467:48:freechips.rocketchip.system.DefaultConfig.fir@220937.4]
  wire  _T_725; // @[Monitor.scala 467:12:freechips.rocketchip.system.DefaultConfig.fir@220939.4]
  wire  _T_726; // @[Monitor.scala 467:12:freechips.rocketchip.system.DefaultConfig.fir@220940.4]
  wire [31:0] _T_728; // @[Monitor.scala 469:26:freechips.rocketchip.system.DefaultConfig.fir@220946.4]
  wire  _T_731; // @[Monitor.scala 470:27:freechips.rocketchip.system.DefaultConfig.fir@220950.4]
  wire  _GEN_19; // @[Monitor.scala 41:14:freechips.rocketchip.system.DefaultConfig.fir@219893.10]
  wire  _GEN_33; // @[Monitor.scala 52:14:freechips.rocketchip.system.DefaultConfig.fir@219965.10]
  wire  _GEN_49; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220048.10]
  wire  _GEN_59; // @[Monitor.scala 73:14:freechips.rocketchip.system.DefaultConfig.fir@220107.10]
  wire  _GEN_67; // @[Monitor.scala 81:14:freechips.rocketchip.system.DefaultConfig.fir@220158.10]
  wire  _GEN_75; // @[Monitor.scala 89:14:freechips.rocketchip.system.DefaultConfig.fir@220208.10]
  wire  _GEN_83; // @[Monitor.scala 97:14:freechips.rocketchip.system.DefaultConfig.fir@220256.10]
  wire  _GEN_91; // @[Monitor.scala 105:14:freechips.rocketchip.system.DefaultConfig.fir@220304.10]
  wire  _GEN_99; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220374.10]
  wire  _GEN_101; // @[Monitor.scala 273:14:freechips.rocketchip.system.DefaultConfig.fir@220415.10]
  wire  _GEN_105; // @[Monitor.scala 283:14:freechips.rocketchip.system.DefaultConfig.fir@220473.10]
  plusarg_reader #(.FORMAT("tilelink_timeout=%d"), .DEFAULT(0)) plusarg_reader ( // @[PlusArg.scala 42:11:freechips.rocketchip.system.DefaultConfig.fir@220930.4]
    .out(plusarg_reader_out)
  );
  assign _T_36 = 13'h3f << io_in_a_bits_size; // @[package.scala 185:77:freechips.rocketchip.system.DefaultConfig.fir@219810.6]
  assign _T_37 = _T_36[5:0]; // @[package.scala 185:82:freechips.rocketchip.system.DefaultConfig.fir@219811.6]
  assign _T_38 = ~ _T_37; // @[package.scala 185:46:freechips.rocketchip.system.DefaultConfig.fir@219812.6]
  assign _GEN_18 = {{27'd0}, _T_38}; // @[Edges.scala 21:16:freechips.rocketchip.system.DefaultConfig.fir@219813.6]
  assign _T_39 = io_in_a_bits_address & _GEN_18; // @[Edges.scala 21:16:freechips.rocketchip.system.DefaultConfig.fir@219813.6]
  assign _T_40 = _T_39 == 33'h0; // @[Edges.scala 21:24:freechips.rocketchip.system.DefaultConfig.fir@219814.6]
  assign _T_42 = io_in_a_bits_size[1:0]; // @[OneHot.scala 51:49:freechips.rocketchip.system.DefaultConfig.fir@219816.6]
  assign _T_43 = 4'h1 << _T_42; // @[OneHot.scala 52:12:freechips.rocketchip.system.DefaultConfig.fir@219817.6]
  assign _T_44 = _T_43[2:0]; // @[OneHot.scala 52:27:freechips.rocketchip.system.DefaultConfig.fir@219818.6]
  assign _T_45 = _T_44 | 3'h1; // @[Misc.scala 206:81:freechips.rocketchip.system.DefaultConfig.fir@219819.6]
  assign _T_46 = io_in_a_bits_size >= 3'h3; // @[Misc.scala 210:21:freechips.rocketchip.system.DefaultConfig.fir@219820.6]
  assign _T_47 = _T_45[2]; // @[Misc.scala 213:26:freechips.rocketchip.system.DefaultConfig.fir@219821.6]
  assign _T_48 = io_in_a_bits_address[2]; // @[Misc.scala 214:26:freechips.rocketchip.system.DefaultConfig.fir@219822.6]
  assign _T_49 = _T_48 == 1'h0; // @[Misc.scala 215:20:freechips.rocketchip.system.DefaultConfig.fir@219823.6]
  assign _T_51 = _T_47 & _T_49; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219825.6]
  assign _T_52 = _T_46 | _T_51; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219826.6]
  assign _T_54 = _T_47 & _T_48; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219828.6]
  assign _T_55 = _T_46 | _T_54; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219829.6]
  assign _T_56 = _T_45[1]; // @[Misc.scala 213:26:freechips.rocketchip.system.DefaultConfig.fir@219830.6]
  assign _T_57 = io_in_a_bits_address[1]; // @[Misc.scala 214:26:freechips.rocketchip.system.DefaultConfig.fir@219831.6]
  assign _T_58 = _T_57 == 1'h0; // @[Misc.scala 215:20:freechips.rocketchip.system.DefaultConfig.fir@219832.6]
  assign _T_59 = _T_49 & _T_58; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219833.6]
  assign _T_60 = _T_56 & _T_59; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219834.6]
  assign _T_61 = _T_52 | _T_60; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219835.6]
  assign _T_62 = _T_49 & _T_57; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219836.6]
  assign _T_63 = _T_56 & _T_62; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219837.6]
  assign _T_64 = _T_52 | _T_63; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219838.6]
  assign _T_65 = _T_48 & _T_58; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219839.6]
  assign _T_66 = _T_56 & _T_65; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219840.6]
  assign _T_67 = _T_55 | _T_66; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219841.6]
  assign _T_68 = _T_48 & _T_57; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219842.6]
  assign _T_69 = _T_56 & _T_68; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219843.6]
  assign _T_70 = _T_55 | _T_69; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219844.6]
  assign _T_71 = _T_45[0]; // @[Misc.scala 213:26:freechips.rocketchip.system.DefaultConfig.fir@219845.6]
  assign _T_72 = io_in_a_bits_address[0]; // @[Misc.scala 214:26:freechips.rocketchip.system.DefaultConfig.fir@219846.6]
  assign _T_73 = _T_72 == 1'h0; // @[Misc.scala 215:20:freechips.rocketchip.system.DefaultConfig.fir@219847.6]
  assign _T_74 = _T_59 & _T_73; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219848.6]
  assign _T_75 = _T_71 & _T_74; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219849.6]
  assign _T_76 = _T_61 | _T_75; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219850.6]
  assign _T_77 = _T_59 & _T_72; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219851.6]
  assign _T_78 = _T_71 & _T_77; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219852.6]
  assign _T_79 = _T_61 | _T_78; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219853.6]
  assign _T_80 = _T_62 & _T_73; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219854.6]
  assign _T_81 = _T_71 & _T_80; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219855.6]
  assign _T_82 = _T_64 | _T_81; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219856.6]
  assign _T_83 = _T_62 & _T_72; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219857.6]
  assign _T_84 = _T_71 & _T_83; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219858.6]
  assign _T_85 = _T_64 | _T_84; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219859.6]
  assign _T_86 = _T_65 & _T_73; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219860.6]
  assign _T_87 = _T_71 & _T_86; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219861.6]
  assign _T_88 = _T_67 | _T_87; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219862.6]
  assign _T_89 = _T_65 & _T_72; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219863.6]
  assign _T_90 = _T_71 & _T_89; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219864.6]
  assign _T_91 = _T_67 | _T_90; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219865.6]
  assign _T_92 = _T_68 & _T_73; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219866.6]
  assign _T_93 = _T_71 & _T_92; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219867.6]
  assign _T_94 = _T_70 | _T_93; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219868.6]
  assign _T_95 = _T_68 & _T_72; // @[Misc.scala 218:27:freechips.rocketchip.system.DefaultConfig.fir@219869.6]
  assign _T_96 = _T_71 & _T_95; // @[Misc.scala 219:38:freechips.rocketchip.system.DefaultConfig.fir@219870.6]
  assign _T_97 = _T_70 | _T_96; // @[Misc.scala 219:29:freechips.rocketchip.system.DefaultConfig.fir@219871.6]
  assign _T_98 = {_T_79,_T_76}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219872.6]
  assign _T_99 = {_T_85,_T_82}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219873.6]
  assign _T_100 = {_T_99,_T_98}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219874.6]
  assign _T_101 = {_T_91,_T_88}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219875.6]
  assign _T_102 = {_T_97,_T_94}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219876.6]
  assign _T_103 = {_T_102,_T_101}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219877.6]
  assign _T_104 = {_T_103,_T_100}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@219878.6]
  assign _T_105 = io_in_a_bits_opcode == 3'h6; // @[Monitor.scala 40:25:freechips.rocketchip.system.DefaultConfig.fir@219879.6]
  assign _T_107 = io_in_a_bits_address ^ 33'h100000000; // @[Parameters.scala 121:31:freechips.rocketchip.system.DefaultConfig.fir@219882.8]
  assign _T_108 = {1'b0,$signed(_T_107)}; // @[Parameters.scala 121:49:freechips.rocketchip.system.DefaultConfig.fir@219883.8]
  assign _T_109 = $signed(_T_108) & $signed(-34'sh10000000); // @[Parameters.scala 121:52:freechips.rocketchip.system.DefaultConfig.fir@219884.8]
  assign _T_110 = $signed(_T_109); // @[Parameters.scala 121:52:freechips.rocketchip.system.DefaultConfig.fir@219885.8]
  assign _T_111 = $signed(_T_110) == $signed(34'sh0); // @[Parameters.scala 121:67:freechips.rocketchip.system.DefaultConfig.fir@219886.8]
  assign _T_116 = reset == 1'h0; // @[Monitor.scala 41:14:freechips.rocketchip.system.DefaultConfig.fir@219891.8]
  assign _T_125 = _T_46 | reset; // @[Monitor.scala 44:14:freechips.rocketchip.system.DefaultConfig.fir@219912.8]
  assign _T_126 = _T_125 == 1'h0; // @[Monitor.scala 44:14:freechips.rocketchip.system.DefaultConfig.fir@219913.8]
  assign _T_128 = _T_40 | reset; // @[Monitor.scala 45:14:freechips.rocketchip.system.DefaultConfig.fir@219919.8]
  assign _T_129 = _T_128 == 1'h0; // @[Monitor.scala 45:14:freechips.rocketchip.system.DefaultConfig.fir@219920.8]
  assign _T_130 = io_in_a_bits_param <= 3'h2; // @[Bundles.scala 109:27:freechips.rocketchip.system.DefaultConfig.fir@219925.8]
  assign _T_132 = _T_130 | reset; // @[Monitor.scala 46:14:freechips.rocketchip.system.DefaultConfig.fir@219927.8]
  assign _T_133 = _T_132 == 1'h0; // @[Monitor.scala 46:14:freechips.rocketchip.system.DefaultConfig.fir@219928.8]
  assign _T_134 = ~ io_in_a_bits_mask; // @[Monitor.scala 47:15:freechips.rocketchip.system.DefaultConfig.fir@219933.8]
  assign _T_135 = _T_134 == 8'h0; // @[Monitor.scala 47:28:freechips.rocketchip.system.DefaultConfig.fir@219934.8]
  assign _T_137 = _T_135 | reset; // @[Monitor.scala 47:14:freechips.rocketchip.system.DefaultConfig.fir@219936.8]
  assign _T_138 = _T_137 == 1'h0; // @[Monitor.scala 47:14:freechips.rocketchip.system.DefaultConfig.fir@219937.8]
  assign _T_139 = io_in_a_bits_corrupt == 1'h0; // @[Monitor.scala 48:15:freechips.rocketchip.system.DefaultConfig.fir@219942.8]
  assign _T_141 = _T_139 | reset; // @[Monitor.scala 48:14:freechips.rocketchip.system.DefaultConfig.fir@219944.8]
  assign _T_142 = _T_141 == 1'h0; // @[Monitor.scala 48:14:freechips.rocketchip.system.DefaultConfig.fir@219945.8]
  assign _T_143 = io_in_a_bits_opcode == 3'h7; // @[Monitor.scala 51:25:freechips.rocketchip.system.DefaultConfig.fir@219951.6]
  assign _T_172 = io_in_a_bits_param != 3'h0; // @[Monitor.scala 58:28:freechips.rocketchip.system.DefaultConfig.fir@220005.8]
  assign _T_174 = _T_172 | reset; // @[Monitor.scala 58:14:freechips.rocketchip.system.DefaultConfig.fir@220007.8]
  assign _T_175 = _T_174 == 1'h0; // @[Monitor.scala 58:14:freechips.rocketchip.system.DefaultConfig.fir@220008.8]
  assign _T_185 = io_in_a_bits_opcode == 3'h4; // @[Monitor.scala 63:25:freechips.rocketchip.system.DefaultConfig.fir@220031.6]
  assign _T_187 = io_in_a_bits_size <= 3'h6; // @[Parameters.scala 90:42:freechips.rocketchip.system.DefaultConfig.fir@220034.8]
  assign _T_195 = _T_187 & _T_111; // @[Parameters.scala 168:56:freechips.rocketchip.system.DefaultConfig.fir@220042.8]
  assign _T_198 = _T_195 | reset; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220045.8]
  assign _T_199 = _T_198 == 1'h0; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220046.8]
  assign _T_206 = io_in_a_bits_param == 3'h0; // @[Monitor.scala 67:28:freechips.rocketchip.system.DefaultConfig.fir@220065.8]
  assign _T_208 = _T_206 | reset; // @[Monitor.scala 67:14:freechips.rocketchip.system.DefaultConfig.fir@220067.8]
  assign _T_209 = _T_208 == 1'h0; // @[Monitor.scala 67:14:freechips.rocketchip.system.DefaultConfig.fir@220068.8]
  assign _T_210 = io_in_a_bits_mask == _T_104; // @[Monitor.scala 68:27:freechips.rocketchip.system.DefaultConfig.fir@220073.8]
  assign _T_212 = _T_210 | reset; // @[Monitor.scala 68:14:freechips.rocketchip.system.DefaultConfig.fir@220075.8]
  assign _T_213 = _T_212 == 1'h0; // @[Monitor.scala 68:14:freechips.rocketchip.system.DefaultConfig.fir@220076.8]
  assign _T_218 = io_in_a_bits_opcode == 3'h0; // @[Monitor.scala 72:25:freechips.rocketchip.system.DefaultConfig.fir@220090.6]
  assign _T_247 = io_in_a_bits_opcode == 3'h1; // @[Monitor.scala 80:25:freechips.rocketchip.system.DefaultConfig.fir@220141.6]
  assign _T_272 = ~ _T_104; // @[Monitor.scala 85:30:freechips.rocketchip.system.DefaultConfig.fir@220183.8]
  assign _T_273 = io_in_a_bits_mask & _T_272; // @[Monitor.scala 85:28:freechips.rocketchip.system.DefaultConfig.fir@220184.8]
  assign _T_274 = _T_273 == 8'h0; // @[Monitor.scala 85:37:freechips.rocketchip.system.DefaultConfig.fir@220185.8]
  assign _T_276 = _T_274 | reset; // @[Monitor.scala 85:14:freechips.rocketchip.system.DefaultConfig.fir@220187.8]
  assign _T_277 = _T_276 == 1'h0; // @[Monitor.scala 85:14:freechips.rocketchip.system.DefaultConfig.fir@220188.8]
  assign _T_278 = io_in_a_bits_opcode == 3'h2; // @[Monitor.scala 88:25:freechips.rocketchip.system.DefaultConfig.fir@220194.6]
  assign _T_296 = io_in_a_bits_param <= 3'h4; // @[Bundles.scala 139:33:freechips.rocketchip.system.DefaultConfig.fir@220225.8]
  assign _T_298 = _T_296 | reset; // @[Monitor.scala 92:14:freechips.rocketchip.system.DefaultConfig.fir@220227.8]
  assign _T_299 = _T_298 == 1'h0; // @[Monitor.scala 92:14:freechips.rocketchip.system.DefaultConfig.fir@220228.8]
  assign _T_304 = io_in_a_bits_opcode == 3'h3; // @[Monitor.scala 96:25:freechips.rocketchip.system.DefaultConfig.fir@220242.6]
  assign _T_322 = io_in_a_bits_param <= 3'h3; // @[Bundles.scala 146:30:freechips.rocketchip.system.DefaultConfig.fir@220273.8]
  assign _T_324 = _T_322 | reset; // @[Monitor.scala 100:14:freechips.rocketchip.system.DefaultConfig.fir@220275.8]
  assign _T_325 = _T_324 == 1'h0; // @[Monitor.scala 100:14:freechips.rocketchip.system.DefaultConfig.fir@220276.8]
  assign _T_330 = io_in_a_bits_opcode == 3'h5; // @[Monitor.scala 104:25:freechips.rocketchip.system.DefaultConfig.fir@220290.6]
  assign _T_356 = io_in_d_bits_opcode <= 3'h6; // @[Bundles.scala 43:24:freechips.rocketchip.system.DefaultConfig.fir@220340.6]
  assign _T_358 = _T_356 | reset; // @[Monitor.scala 256:12:freechips.rocketchip.system.DefaultConfig.fir@220342.6]
  assign _T_359 = _T_358 == 1'h0; // @[Monitor.scala 256:12:freechips.rocketchip.system.DefaultConfig.fir@220343.6]
  assign _T_376 = io_in_d_bits_opcode == 3'h6; // @[Monitor.scala 263:25:freechips.rocketchip.system.DefaultConfig.fir@220360.6]
  assign _T_380 = io_in_d_bits_size >= 3'h3; // @[Monitor.scala 265:27:freechips.rocketchip.system.DefaultConfig.fir@220369.8]
  assign _T_382 = _T_380 | reset; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220371.8]
  assign _T_383 = _T_382 == 1'h0; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220372.8]
  assign _T_396 = io_in_d_bits_opcode == 3'h4; // @[Monitor.scala 271:25:freechips.rocketchip.system.DefaultConfig.fir@220402.6]
  assign _T_424 = io_in_d_bits_opcode == 3'h5; // @[Monitor.scala 281:25:freechips.rocketchip.system.DefaultConfig.fir@220460.6]
  assign _T_517 = io_in_a_ready & io_in_a_valid; // @[Bundles.scala 283:22:freechips.rocketchip.system.DefaultConfig.fir@220650.4]
  assign _T_522 = _T_38[5:3]; // @[Edges.scala 220:59:freechips.rocketchip.system.DefaultConfig.fir@220655.4]
  assign _T_523 = io_in_a_bits_opcode[2]; // @[Edges.scala 92:37:freechips.rocketchip.system.DefaultConfig.fir@220656.4]
  assign _T_524 = _T_523 == 1'h0; // @[Edges.scala 92:28:freechips.rocketchip.system.DefaultConfig.fir@220657.4]
  assign _T_528 = _T_527 - 3'h1; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220660.4]
  assign _T_529 = $unsigned(_T_528); // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220661.4]
  assign _T_530 = _T_529[2:0]; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220662.4]
  assign _T_531 = _T_527 == 3'h0; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220663.4]
  assign _T_549 = _T_531 == 1'h0; // @[Monitor.scala 342:22:freechips.rocketchip.system.DefaultConfig.fir@220679.4]
  assign _T_550 = io_in_a_valid & _T_549; // @[Monitor.scala 342:19:freechips.rocketchip.system.DefaultConfig.fir@220680.4]
  assign _T_551 = io_in_a_bits_opcode == _T_540; // @[Monitor.scala 343:29:freechips.rocketchip.system.DefaultConfig.fir@220682.6]
  assign _T_553 = _T_551 | reset; // @[Monitor.scala 343:14:freechips.rocketchip.system.DefaultConfig.fir@220684.6]
  assign _T_554 = _T_553 == 1'h0; // @[Monitor.scala 343:14:freechips.rocketchip.system.DefaultConfig.fir@220685.6]
  assign _T_555 = io_in_a_bits_param == _T_542; // @[Monitor.scala 344:29:freechips.rocketchip.system.DefaultConfig.fir@220690.6]
  assign _T_557 = _T_555 | reset; // @[Monitor.scala 344:14:freechips.rocketchip.system.DefaultConfig.fir@220692.6]
  assign _T_558 = _T_557 == 1'h0; // @[Monitor.scala 344:14:freechips.rocketchip.system.DefaultConfig.fir@220693.6]
  assign _T_559 = io_in_a_bits_size == _T_544; // @[Monitor.scala 345:29:freechips.rocketchip.system.DefaultConfig.fir@220698.6]
  assign _T_561 = _T_559 | reset; // @[Monitor.scala 345:14:freechips.rocketchip.system.DefaultConfig.fir@220700.6]
  assign _T_562 = _T_561 == 1'h0; // @[Monitor.scala 345:14:freechips.rocketchip.system.DefaultConfig.fir@220701.6]
  assign _T_563 = io_in_a_bits_source == _T_546; // @[Monitor.scala 346:29:freechips.rocketchip.system.DefaultConfig.fir@220706.6]
  assign _T_565 = _T_563 | reset; // @[Monitor.scala 346:14:freechips.rocketchip.system.DefaultConfig.fir@220708.6]
  assign _T_566 = _T_565 == 1'h0; // @[Monitor.scala 346:14:freechips.rocketchip.system.DefaultConfig.fir@220709.6]
  assign _T_567 = io_in_a_bits_address == _T_548; // @[Monitor.scala 347:29:freechips.rocketchip.system.DefaultConfig.fir@220714.6]
  assign _T_569 = _T_567 | reset; // @[Monitor.scala 347:14:freechips.rocketchip.system.DefaultConfig.fir@220716.6]
  assign _T_570 = _T_569 == 1'h0; // @[Monitor.scala 347:14:freechips.rocketchip.system.DefaultConfig.fir@220717.6]
  assign _T_572 = _T_517 & _T_531; // @[Monitor.scala 349:20:freechips.rocketchip.system.DefaultConfig.fir@220724.4]
  assign _T_573 = io_in_d_ready & io_in_d_valid; // @[Bundles.scala 283:22:freechips.rocketchip.system.DefaultConfig.fir@220732.4]
  assign _T_575 = 13'h3f << io_in_d_bits_size; // @[package.scala 185:77:freechips.rocketchip.system.DefaultConfig.fir@220734.4]
  assign _T_576 = _T_575[5:0]; // @[package.scala 185:82:freechips.rocketchip.system.DefaultConfig.fir@220735.4]
  assign _T_577 = ~ _T_576; // @[package.scala 185:46:freechips.rocketchip.system.DefaultConfig.fir@220736.4]
  assign _T_578 = _T_577[5:3]; // @[Edges.scala 220:59:freechips.rocketchip.system.DefaultConfig.fir@220737.4]
  assign _T_579 = io_in_d_bits_opcode[0]; // @[Edges.scala 106:36:freechips.rocketchip.system.DefaultConfig.fir@220738.4]
  assign _T_583 = _T_582 - 3'h1; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220741.4]
  assign _T_584 = $unsigned(_T_583); // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220742.4]
  assign _T_585 = _T_584[2:0]; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220743.4]
  assign _T_586 = _T_582 == 3'h0; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220744.4]
  assign _T_606 = _T_586 == 1'h0; // @[Monitor.scala 412:22:freechips.rocketchip.system.DefaultConfig.fir@220761.4]
  assign _T_607 = io_in_d_valid & _T_606; // @[Monitor.scala 412:19:freechips.rocketchip.system.DefaultConfig.fir@220762.4]
  assign _T_608 = io_in_d_bits_opcode == _T_595; // @[Monitor.scala 413:29:freechips.rocketchip.system.DefaultConfig.fir@220764.6]
  assign _T_610 = _T_608 | reset; // @[Monitor.scala 413:14:freechips.rocketchip.system.DefaultConfig.fir@220766.6]
  assign _T_611 = _T_610 == 1'h0; // @[Monitor.scala 413:14:freechips.rocketchip.system.DefaultConfig.fir@220767.6]
  assign _T_616 = io_in_d_bits_size == _T_599; // @[Monitor.scala 415:29:freechips.rocketchip.system.DefaultConfig.fir@220780.6]
  assign _T_618 = _T_616 | reset; // @[Monitor.scala 415:14:freechips.rocketchip.system.DefaultConfig.fir@220782.6]
  assign _T_619 = _T_618 == 1'h0; // @[Monitor.scala 415:14:freechips.rocketchip.system.DefaultConfig.fir@220783.6]
  assign _T_620 = io_in_d_bits_source == _T_601; // @[Monitor.scala 416:29:freechips.rocketchip.system.DefaultConfig.fir@220788.6]
  assign _T_622 = _T_620 | reset; // @[Monitor.scala 416:14:freechips.rocketchip.system.DefaultConfig.fir@220790.6]
  assign _T_623 = _T_622 == 1'h0; // @[Monitor.scala 416:14:freechips.rocketchip.system.DefaultConfig.fir@220791.6]
  assign _T_633 = _T_573 & _T_586; // @[Monitor.scala 420:20:freechips.rocketchip.system.DefaultConfig.fir@220814.4]
  assign _T_647 = _T_646 - 3'h1; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220834.4]
  assign _T_648 = $unsigned(_T_647); // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220835.4]
  assign _T_649 = _T_648[2:0]; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220836.4]
  assign _T_650 = _T_646 == 3'h0; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220837.4]
  assign _T_668 = _T_667 - 3'h1; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220857.4]
  assign _T_669 = $unsigned(_T_668); // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220858.4]
  assign _T_670 = _T_669[2:0]; // @[Edges.scala 230:28:freechips.rocketchip.system.DefaultConfig.fir@220859.4]
  assign _T_671 = _T_667 == 3'h0; // @[Edges.scala 231:25:freechips.rocketchip.system.DefaultConfig.fir@220860.4]
  assign _T_682 = _T_517 & _T_650; // @[Monitor.scala 446:27:freechips.rocketchip.system.DefaultConfig.fir@220875.4]
  assign _T_684 = 64'h1 << io_in_a_bits_source; // @[OneHot.scala 45:35:freechips.rocketchip.system.DefaultConfig.fir@220878.6]
  assign _T_685 = _T_635 >> io_in_a_bits_source; // @[Monitor.scala 448:23:freechips.rocketchip.system.DefaultConfig.fir@220880.6]
  assign _T_686 = _T_685[0]; // @[Monitor.scala 448:23:freechips.rocketchip.system.DefaultConfig.fir@220881.6]
  assign _T_687 = _T_686 == 1'h0; // @[Monitor.scala 448:14:freechips.rocketchip.system.DefaultConfig.fir@220882.6]
  assign _T_689 = _T_687 | reset; // @[Monitor.scala 448:13:freechips.rocketchip.system.DefaultConfig.fir@220884.6]
  assign _T_690 = _T_689 == 1'h0; // @[Monitor.scala 448:13:freechips.rocketchip.system.DefaultConfig.fir@220885.6]
  assign _GEN_15 = _T_682 ? _T_684 : 64'h0; // @[Monitor.scala 446:72:freechips.rocketchip.system.DefaultConfig.fir@220877.4]
  assign _T_695 = _T_573 & _T_671; // @[Monitor.scala 453:27:freechips.rocketchip.system.DefaultConfig.fir@220896.4]
  assign _T_697 = _T_376 == 1'h0; // @[Monitor.scala 453:75:freechips.rocketchip.system.DefaultConfig.fir@220898.4]
  assign _T_698 = _T_695 & _T_697; // @[Monitor.scala 453:72:freechips.rocketchip.system.DefaultConfig.fir@220899.4]
  assign _T_699 = 64'h1 << io_in_d_bits_source; // @[OneHot.scala 45:35:freechips.rocketchip.system.DefaultConfig.fir@220901.6]
  assign _T_700 = _GEN_15 | _T_635; // @[Monitor.scala 455:21:freechips.rocketchip.system.DefaultConfig.fir@220903.6]
  assign _T_701 = _T_700 >> io_in_d_bits_source; // @[Monitor.scala 455:32:freechips.rocketchip.system.DefaultConfig.fir@220904.6]
  assign _T_702 = _T_701[0]; // @[Monitor.scala 455:32:freechips.rocketchip.system.DefaultConfig.fir@220905.6]
  assign _T_704 = _T_702 | reset; // @[Monitor.scala 455:13:freechips.rocketchip.system.DefaultConfig.fir@220907.6]
  assign _T_705 = _T_704 == 1'h0; // @[Monitor.scala 455:13:freechips.rocketchip.system.DefaultConfig.fir@220908.6]
  assign _GEN_16 = _T_698 ? _T_699 : 64'h0; // @[Monitor.scala 453:91:freechips.rocketchip.system.DefaultConfig.fir@220900.4]
  assign _T_706 = _GEN_15 != _GEN_16; // @[Monitor.scala 459:20:freechips.rocketchip.system.DefaultConfig.fir@220914.4]
  assign _T_707 = _GEN_15 != 64'h0; // @[Monitor.scala 459:40:freechips.rocketchip.system.DefaultConfig.fir@220915.4]
  assign _T_708 = _T_707 == 1'h0; // @[Monitor.scala 459:33:freechips.rocketchip.system.DefaultConfig.fir@220916.4]
  assign _T_709 = _T_706 | _T_708; // @[Monitor.scala 459:30:freechips.rocketchip.system.DefaultConfig.fir@220917.4]
  assign _T_711 = _T_709 | reset; // @[Monitor.scala 459:13:freechips.rocketchip.system.DefaultConfig.fir@220919.4]
  assign _T_712 = _T_711 == 1'h0; // @[Monitor.scala 459:13:freechips.rocketchip.system.DefaultConfig.fir@220920.4]
  assign _T_713 = _T_635 | _GEN_15; // @[Monitor.scala 462:27:freechips.rocketchip.system.DefaultConfig.fir@220925.4]
  assign _T_714 = ~ _GEN_16; // @[Monitor.scala 462:38:freechips.rocketchip.system.DefaultConfig.fir@220926.4]
  assign _T_715 = _T_713 & _T_714; // @[Monitor.scala 462:36:freechips.rocketchip.system.DefaultConfig.fir@220927.4]
  assign _T_718 = _T_635 != 64'h0; // @[Monitor.scala 467:23:freechips.rocketchip.system.DefaultConfig.fir@220932.4]
  assign _T_719 = _T_718 == 1'h0; // @[Monitor.scala 467:13:freechips.rocketchip.system.DefaultConfig.fir@220933.4]
  assign _T_720 = plusarg_reader_out == 32'h0; // @[Monitor.scala 467:36:freechips.rocketchip.system.DefaultConfig.fir@220934.4]
  assign _T_721 = _T_719 | _T_720; // @[Monitor.scala 467:27:freechips.rocketchip.system.DefaultConfig.fir@220935.4]
  assign _T_722 = _T_717 < plusarg_reader_out; // @[Monitor.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@220936.4]
  assign _T_723 = _T_721 | _T_722; // @[Monitor.scala 467:48:freechips.rocketchip.system.DefaultConfig.fir@220937.4]
  assign _T_725 = _T_723 | reset; // @[Monitor.scala 467:12:freechips.rocketchip.system.DefaultConfig.fir@220939.4]
  assign _T_726 = _T_725 == 1'h0; // @[Monitor.scala 467:12:freechips.rocketchip.system.DefaultConfig.fir@220940.4]
  assign _T_728 = _T_717 + 32'h1; // @[Monitor.scala 469:26:freechips.rocketchip.system.DefaultConfig.fir@220946.4]
  assign _T_731 = _T_517 | _T_573; // @[Monitor.scala 470:27:freechips.rocketchip.system.DefaultConfig.fir@220950.4]
  assign _GEN_19 = io_in_a_valid & _T_105; // @[Monitor.scala 41:14:freechips.rocketchip.system.DefaultConfig.fir@219893.10]
  assign _GEN_33 = io_in_a_valid & _T_143; // @[Monitor.scala 52:14:freechips.rocketchip.system.DefaultConfig.fir@219965.10]
  assign _GEN_49 = io_in_a_valid & _T_185; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220048.10]
  assign _GEN_59 = io_in_a_valid & _T_218; // @[Monitor.scala 73:14:freechips.rocketchip.system.DefaultConfig.fir@220107.10]
  assign _GEN_67 = io_in_a_valid & _T_247; // @[Monitor.scala 81:14:freechips.rocketchip.system.DefaultConfig.fir@220158.10]
  assign _GEN_75 = io_in_a_valid & _T_278; // @[Monitor.scala 89:14:freechips.rocketchip.system.DefaultConfig.fir@220208.10]
  assign _GEN_83 = io_in_a_valid & _T_304; // @[Monitor.scala 97:14:freechips.rocketchip.system.DefaultConfig.fir@220256.10]
  assign _GEN_91 = io_in_a_valid & _T_330; // @[Monitor.scala 105:14:freechips.rocketchip.system.DefaultConfig.fir@220304.10]
  assign _GEN_99 = io_in_d_valid & _T_376; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220374.10]
  assign _GEN_101 = io_in_d_valid & _T_396; // @[Monitor.scala 273:14:freechips.rocketchip.system.DefaultConfig.fir@220415.10]
  assign _GEN_105 = io_in_d_valid & _T_424; // @[Monitor.scala 283:14:freechips.rocketchip.system.DefaultConfig.fir@220473.10]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_527 = _RAND_0[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_540 = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_542 = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_544 = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_546 = _RAND_4[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {2{`RANDOM}};
  _T_548 = _RAND_5[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_582 = _RAND_6[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_595 = _RAND_7[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_599 = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_601 = _RAND_9[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {2{`RANDOM}};
  _T_635 = _RAND_10[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_646 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_667 = _RAND_12[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  _T_717 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_527 <= 3'h0;
    end else begin
      if (_T_517) begin
        if (_T_531) begin
          if (_T_524) begin
            _T_527 <= _T_522;
          end else begin
            _T_527 <= 3'h0;
          end
        end else begin
          _T_527 <= _T_530;
        end
      end
    end
    if (_T_572) begin
      _T_540 <= io_in_a_bits_opcode;
    end
    if (_T_572) begin
      _T_542 <= io_in_a_bits_param;
    end
    if (_T_572) begin
      _T_544 <= io_in_a_bits_size;
    end
    if (_T_572) begin
      _T_546 <= io_in_a_bits_source;
    end
    if (_T_572) begin
      _T_548 <= io_in_a_bits_address;
    end
    if (reset) begin
      _T_582 <= 3'h0;
    end else begin
      if (_T_573) begin
        if (_T_586) begin
          if (_T_579) begin
            _T_582 <= _T_578;
          end else begin
            _T_582 <= 3'h0;
          end
        end else begin
          _T_582 <= _T_585;
        end
      end
    end
    if (_T_633) begin
      _T_595 <= io_in_d_bits_opcode;
    end
    if (_T_633) begin
      _T_599 <= io_in_d_bits_size;
    end
    if (_T_633) begin
      _T_601 <= io_in_d_bits_source;
    end
    if (reset) begin
      _T_635 <= 64'h0;
    end else begin
      _T_635 <= _T_715;
    end
    if (reset) begin
      _T_646 <= 3'h0;
    end else begin
      if (_T_517) begin
        if (_T_650) begin
          if (_T_524) begin
            _T_646 <= _T_522;
          end else begin
            _T_646 <= 3'h0;
          end
        end else begin
          _T_646 <= _T_649;
        end
      end
    end
    if (reset) begin
      _T_667 <= 3'h0;
    end else begin
      if (_T_573) begin
        if (_T_671) begin
          if (_T_579) begin
            _T_667 <= _T_578;
          end else begin
            _T_667 <= 3'h0;
          end
        end else begin
          _T_667 <= _T_670;
        end
      end
    end
    if (reset) begin
      _T_717 <= 32'h0;
    end else begin
      if (_T_731) begin
        _T_717 <= 32'h0;
      end else begin
        _T_717 <= _T_728;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel has invalid opcode (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:33 assert (TLMessages.isA(bundle.opcode), \"'A' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 33:12:freechips.rocketchip.system.DefaultConfig.fir@219795.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 33:12:freechips.rocketchip.system.DefaultConfig.fir@219796.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:41 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquireBlock type unsupported by manager\" + extra)\n"); // @[Monitor.scala 41:14:freechips.rocketchip.system.DefaultConfig.fir@219893.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fatal; // @[Monitor.scala 41:14:freechips.rocketchip.system.DefaultConfig.fir@219894.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquireBlock from a client which does not support Probe (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:42 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquireBlock from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 42:14:freechips.rocketchip.system.DefaultConfig.fir@219900.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_116) begin
          $fatal; // @[Monitor.scala 42:14:freechips.rocketchip.system.DefaultConfig.fir@219901.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:43 assert (source_ok, \"'A' channel AcquireBlock carries invalid source ID\" + extra)\n"); // @[Monitor.scala 43:14:freechips.rocketchip.system.DefaultConfig.fir@219907.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 43:14:freechips.rocketchip.system.DefaultConfig.fir@219908.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_126) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock smaller than a beat (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:44 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquireBlock smaller than a beat\" + extra)\n"); // @[Monitor.scala 44:14:freechips.rocketchip.system.DefaultConfig.fir@219915.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_126) begin
          $fatal; // @[Monitor.scala 44:14:freechips.rocketchip.system.DefaultConfig.fir@219916.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:45 assert (is_aligned, \"'A' channel AcquireBlock address not aligned to size\" + extra)\n"); // @[Monitor.scala 45:14:freechips.rocketchip.system.DefaultConfig.fir@219922.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_129) begin
          $fatal; // @[Monitor.scala 45:14:freechips.rocketchip.system.DefaultConfig.fir@219923.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock carries invalid grow param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:46 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquireBlock carries invalid grow param\" + extra)\n"); // @[Monitor.scala 46:14:freechips.rocketchip.system.DefaultConfig.fir@219930.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_133) begin
          $fatal; // @[Monitor.scala 46:14:freechips.rocketchip.system.DefaultConfig.fir@219931.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_138) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:47 assert (~bundle.mask === UInt(0), \"'A' channel AcquireBlock contains invalid mask\" + extra)\n"); // @[Monitor.scala 47:14:freechips.rocketchip.system.DefaultConfig.fir@219939.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_138) begin
          $fatal; // @[Monitor.scala 47:14:freechips.rocketchip.system.DefaultConfig.fir@219940.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_19 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquireBlock is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:48 assert (!bundle.corrupt, \"'A' channel AcquireBlock is corrupt\" + extra)\n"); // @[Monitor.scala 48:14:freechips.rocketchip.system.DefaultConfig.fir@219947.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_19 & _T_142) begin
          $fatal; // @[Monitor.scala 48:14:freechips.rocketchip.system.DefaultConfig.fir@219948.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:52 assert (edge.manager.supportsAcquireBSafe(edge.address(bundle), bundle.size), \"'A' channel carries AcquirePerm type unsupported by manager\" + extra)\n"); // @[Monitor.scala 52:14:freechips.rocketchip.system.DefaultConfig.fir@219965.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_116) begin
          $fatal; // @[Monitor.scala 52:14:freechips.rocketchip.system.DefaultConfig.fir@219966.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries AcquirePerm from a client which does not support Probe (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:53 assert (edge.client.supportsProbe(edge.source(bundle), bundle.size), \"'A' channel carries AcquirePerm from a client which does not support Probe\" + extra)\n"); // @[Monitor.scala 53:14:freechips.rocketchip.system.DefaultConfig.fir@219972.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_116) begin
          $fatal; // @[Monitor.scala 53:14:freechips.rocketchip.system.DefaultConfig.fir@219973.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:54 assert (source_ok, \"'A' channel AcquirePerm carries invalid source ID\" + extra)\n"); // @[Monitor.scala 54:14:freechips.rocketchip.system.DefaultConfig.fir@219979.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 54:14:freechips.rocketchip.system.DefaultConfig.fir@219980.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_126) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm smaller than a beat (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:55 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'A' channel AcquirePerm smaller than a beat\" + extra)\n"); // @[Monitor.scala 55:14:freechips.rocketchip.system.DefaultConfig.fir@219987.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_126) begin
          $fatal; // @[Monitor.scala 55:14:freechips.rocketchip.system.DefaultConfig.fir@219988.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:56 assert (is_aligned, \"'A' channel AcquirePerm address not aligned to size\" + extra)\n"); // @[Monitor.scala 56:14:freechips.rocketchip.system.DefaultConfig.fir@219994.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_129) begin
          $fatal; // @[Monitor.scala 56:14:freechips.rocketchip.system.DefaultConfig.fir@219995.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_133) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm carries invalid grow param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:57 assert (TLPermissions.isGrow(bundle.param), \"'A' channel AcquirePerm carries invalid grow param\" + extra)\n"); // @[Monitor.scala 57:14:freechips.rocketchip.system.DefaultConfig.fir@220002.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_133) begin
          $fatal; // @[Monitor.scala 57:14:freechips.rocketchip.system.DefaultConfig.fir@220003.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_175) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm requests NtoB (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:58 assert (bundle.param =/= TLPermissions.NtoB, \"'A' channel AcquirePerm requests NtoB\" + extra)\n"); // @[Monitor.scala 58:14:freechips.rocketchip.system.DefaultConfig.fir@220010.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_175) begin
          $fatal; // @[Monitor.scala 58:14:freechips.rocketchip.system.DefaultConfig.fir@220011.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_138) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:59 assert (~bundle.mask === UInt(0), \"'A' channel AcquirePerm contains invalid mask\" + extra)\n"); // @[Monitor.scala 59:14:freechips.rocketchip.system.DefaultConfig.fir@220019.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_138) begin
          $fatal; // @[Monitor.scala 59:14:freechips.rocketchip.system.DefaultConfig.fir@220020.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_33 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel AcquirePerm is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:60 assert (!bundle.corrupt, \"'A' channel AcquirePerm is corrupt\" + extra)\n"); // @[Monitor.scala 60:14:freechips.rocketchip.system.DefaultConfig.fir@220027.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_33 & _T_142) begin
          $fatal; // @[Monitor.scala 60:14:freechips.rocketchip.system.DefaultConfig.fir@220028.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_199) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Get type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:64 assert (edge.manager.supportsGetSafe(edge.address(bundle), bundle.size), \"'A' channel carries Get type unsupported by manager\" + extra)\n"); // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220048.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_199) begin
          $fatal; // @[Monitor.scala 64:14:freechips.rocketchip.system.DefaultConfig.fir@220049.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:65 assert (source_ok, \"'A' channel Get carries invalid source ID\" + extra)\n"); // @[Monitor.scala 65:14:freechips.rocketchip.system.DefaultConfig.fir@220055.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 65:14:freechips.rocketchip.system.DefaultConfig.fir@220056.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:66 assert (is_aligned, \"'A' channel Get address not aligned to size\" + extra)\n"); // @[Monitor.scala 66:14:freechips.rocketchip.system.DefaultConfig.fir@220062.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_129) begin
          $fatal; // @[Monitor.scala 66:14:freechips.rocketchip.system.DefaultConfig.fir@220063.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_209) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:67 assert (bundle.param === UInt(0), \"'A' channel Get carries invalid param\" + extra)\n"); // @[Monitor.scala 67:14:freechips.rocketchip.system.DefaultConfig.fir@220070.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_209) begin
          $fatal; // @[Monitor.scala 67:14:freechips.rocketchip.system.DefaultConfig.fir@220071.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_213) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:68 assert (bundle.mask === mask, \"'A' channel Get contains invalid mask\" + extra)\n"); // @[Monitor.scala 68:14:freechips.rocketchip.system.DefaultConfig.fir@220078.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_213) begin
          $fatal; // @[Monitor.scala 68:14:freechips.rocketchip.system.DefaultConfig.fir@220079.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_49 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Get is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:69 assert (!bundle.corrupt, \"'A' channel Get is corrupt\" + extra)\n"); // @[Monitor.scala 69:14:freechips.rocketchip.system.DefaultConfig.fir@220086.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_49 & _T_142) begin
          $fatal; // @[Monitor.scala 69:14:freechips.rocketchip.system.DefaultConfig.fir@220087.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_59 & _T_199) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutFull type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:73 assert (edge.manager.supportsPutFullSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutFull type unsupported by manager\" + extra)\n"); // @[Monitor.scala 73:14:freechips.rocketchip.system.DefaultConfig.fir@220107.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_59 & _T_199) begin
          $fatal; // @[Monitor.scala 73:14:freechips.rocketchip.system.DefaultConfig.fir@220108.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:74 assert (source_ok, \"'A' channel PutFull carries invalid source ID\" + extra)\n"); // @[Monitor.scala 74:14:freechips.rocketchip.system.DefaultConfig.fir@220114.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 74:14:freechips.rocketchip.system.DefaultConfig.fir@220115.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_59 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:75 assert (is_aligned, \"'A' channel PutFull address not aligned to size\" + extra)\n"); // @[Monitor.scala 75:14:freechips.rocketchip.system.DefaultConfig.fir@220121.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_59 & _T_129) begin
          $fatal; // @[Monitor.scala 75:14:freechips.rocketchip.system.DefaultConfig.fir@220122.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_59 & _T_209) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:76 assert (bundle.param === UInt(0), \"'A' channel PutFull carries invalid param\" + extra)\n"); // @[Monitor.scala 76:14:freechips.rocketchip.system.DefaultConfig.fir@220129.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_59 & _T_209) begin
          $fatal; // @[Monitor.scala 76:14:freechips.rocketchip.system.DefaultConfig.fir@220130.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_59 & _T_213) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutFull contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:77 assert (bundle.mask === mask, \"'A' channel PutFull contains invalid mask\" + extra)\n"); // @[Monitor.scala 77:14:freechips.rocketchip.system.DefaultConfig.fir@220137.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_59 & _T_213) begin
          $fatal; // @[Monitor.scala 77:14:freechips.rocketchip.system.DefaultConfig.fir@220138.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_199) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries PutPartial type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:81 assert (edge.manager.supportsPutPartialSafe(edge.address(bundle), bundle.size), \"'A' channel carries PutPartial type unsupported by manager\" + extra)\n"); // @[Monitor.scala 81:14:freechips.rocketchip.system.DefaultConfig.fir@220158.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_199) begin
          $fatal; // @[Monitor.scala 81:14:freechips.rocketchip.system.DefaultConfig.fir@220159.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:82 assert (source_ok, \"'A' channel PutPartial carries invalid source ID\" + extra)\n"); // @[Monitor.scala 82:14:freechips.rocketchip.system.DefaultConfig.fir@220165.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 82:14:freechips.rocketchip.system.DefaultConfig.fir@220166.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:83 assert (is_aligned, \"'A' channel PutPartial address not aligned to size\" + extra)\n"); // @[Monitor.scala 83:14:freechips.rocketchip.system.DefaultConfig.fir@220172.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_129) begin
          $fatal; // @[Monitor.scala 83:14:freechips.rocketchip.system.DefaultConfig.fir@220173.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_209) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:84 assert (bundle.param === UInt(0), \"'A' channel PutPartial carries invalid param\" + extra)\n"); // @[Monitor.scala 84:14:freechips.rocketchip.system.DefaultConfig.fir@220180.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_209) begin
          $fatal; // @[Monitor.scala 84:14:freechips.rocketchip.system.DefaultConfig.fir@220181.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_67 & _T_277) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel PutPartial contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:85 assert ((bundle.mask & ~mask) === UInt(0), \"'A' channel PutPartial contains invalid mask\" + extra)\n"); // @[Monitor.scala 85:14:freechips.rocketchip.system.DefaultConfig.fir@220190.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_67 & _T_277) begin
          $fatal; // @[Monitor.scala 85:14:freechips.rocketchip.system.DefaultConfig.fir@220191.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Arithmetic type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:89 assert (edge.manager.supportsArithmeticSafe(edge.address(bundle), bundle.size), \"'A' channel carries Arithmetic type unsupported by manager\" + extra)\n"); // @[Monitor.scala 89:14:freechips.rocketchip.system.DefaultConfig.fir@220208.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_116) begin
          $fatal; // @[Monitor.scala 89:14:freechips.rocketchip.system.DefaultConfig.fir@220209.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:90 assert (source_ok, \"'A' channel Arithmetic carries invalid source ID\" + extra)\n"); // @[Monitor.scala 90:14:freechips.rocketchip.system.DefaultConfig.fir@220215.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 90:14:freechips.rocketchip.system.DefaultConfig.fir@220216.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:91 assert (is_aligned, \"'A' channel Arithmetic address not aligned to size\" + extra)\n"); // @[Monitor.scala 91:14:freechips.rocketchip.system.DefaultConfig.fir@220222.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_129) begin
          $fatal; // @[Monitor.scala 91:14:freechips.rocketchip.system.DefaultConfig.fir@220223.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_299) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic carries invalid opcode param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:92 assert (TLAtomics.isArithmetic(bundle.param), \"'A' channel Arithmetic carries invalid opcode param\" + extra)\n"); // @[Monitor.scala 92:14:freechips.rocketchip.system.DefaultConfig.fir@220230.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_299) begin
          $fatal; // @[Monitor.scala 92:14:freechips.rocketchip.system.DefaultConfig.fir@220231.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_75 & _T_213) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Arithmetic contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:93 assert (bundle.mask === mask, \"'A' channel Arithmetic contains invalid mask\" + extra)\n"); // @[Monitor.scala 93:14:freechips.rocketchip.system.DefaultConfig.fir@220238.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_75 & _T_213) begin
          $fatal; // @[Monitor.scala 93:14:freechips.rocketchip.system.DefaultConfig.fir@220239.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Logical type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:97 assert (edge.manager.supportsLogicalSafe(edge.address(bundle), bundle.size), \"'A' channel carries Logical type unsupported by manager\" + extra)\n"); // @[Monitor.scala 97:14:freechips.rocketchip.system.DefaultConfig.fir@220256.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & _T_116) begin
          $fatal; // @[Monitor.scala 97:14:freechips.rocketchip.system.DefaultConfig.fir@220257.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:98 assert (source_ok, \"'A' channel Logical carries invalid source ID\" + extra)\n"); // @[Monitor.scala 98:14:freechips.rocketchip.system.DefaultConfig.fir@220263.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 98:14:freechips.rocketchip.system.DefaultConfig.fir@220264.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:99 assert (is_aligned, \"'A' channel Logical address not aligned to size\" + extra)\n"); // @[Monitor.scala 99:14:freechips.rocketchip.system.DefaultConfig.fir@220270.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & _T_129) begin
          $fatal; // @[Monitor.scala 99:14:freechips.rocketchip.system.DefaultConfig.fir@220271.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & _T_325) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical carries invalid opcode param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:100 assert (TLAtomics.isLogical(bundle.param), \"'A' channel Logical carries invalid opcode param\" + extra)\n"); // @[Monitor.scala 100:14:freechips.rocketchip.system.DefaultConfig.fir@220278.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & _T_325) begin
          $fatal; // @[Monitor.scala 100:14:freechips.rocketchip.system.DefaultConfig.fir@220279.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_83 & _T_213) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Logical contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:101 assert (bundle.mask === mask, \"'A' channel Logical contains invalid mask\" + extra)\n"); // @[Monitor.scala 101:14:freechips.rocketchip.system.DefaultConfig.fir@220286.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_83 & _T_213) begin
          $fatal; // @[Monitor.scala 101:14:freechips.rocketchip.system.DefaultConfig.fir@220287.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel carries Hint type unsupported by manager (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:105 assert (edge.manager.supportsHintSafe(edge.address(bundle), bundle.size), \"'A' channel carries Hint type unsupported by manager\" + extra)\n"); // @[Monitor.scala 105:14:freechips.rocketchip.system.DefaultConfig.fir@220304.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_116) begin
          $fatal; // @[Monitor.scala 105:14:freechips.rocketchip.system.DefaultConfig.fir@220305.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:106 assert (source_ok, \"'A' channel Hint carries invalid source ID\" + extra)\n"); // @[Monitor.scala 106:14:freechips.rocketchip.system.DefaultConfig.fir@220311.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 106:14:freechips.rocketchip.system.DefaultConfig.fir@220312.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_129) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint address not aligned to size (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:107 assert (is_aligned, \"'A' channel Hint address not aligned to size\" + extra)\n"); // @[Monitor.scala 107:14:freechips.rocketchip.system.DefaultConfig.fir@220318.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_129) begin
          $fatal; // @[Monitor.scala 107:14:freechips.rocketchip.system.DefaultConfig.fir@220319.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_213) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint contains invalid mask (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:108 assert (bundle.mask === mask, \"'A' channel Hint contains invalid mask\" + extra)\n"); // @[Monitor.scala 108:14:freechips.rocketchip.system.DefaultConfig.fir@220326.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_213) begin
          $fatal; // @[Monitor.scala 108:14:freechips.rocketchip.system.DefaultConfig.fir@220327.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_91 & _T_142) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel Hint is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:109 assert (!bundle.corrupt, \"'A' channel Hint is corrupt\" + extra)\n"); // @[Monitor.scala 109:14:freechips.rocketchip.system.DefaultConfig.fir@220334.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_91 & _T_142) begin
          $fatal; // @[Monitor.scala 109:14:freechips.rocketchip.system.DefaultConfig.fir@220335.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_in_d_valid & _T_359) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel has invalid opcode (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:256 assert (TLMessages.isD(bundle.opcode), \"'D' channel has invalid opcode\" + extra)\n"); // @[Monitor.scala 256:12:freechips.rocketchip.system.DefaultConfig.fir@220345.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (io_in_d_valid & _T_359) begin
          $fatal; // @[Monitor.scala 256:12:freechips.rocketchip.system.DefaultConfig.fir@220346.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:264 assert (source_ok, \"'D' channel ReleaseAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 264:14:freechips.rocketchip.system.DefaultConfig.fir@220366.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 264:14:freechips.rocketchip.system.DefaultConfig.fir@220367.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_99 & _T_383) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck smaller than a beat (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:265 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel ReleaseAck smaller than a beat\" + extra)\n"); // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220374.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_99 & _T_383) begin
          $fatal; // @[Monitor.scala 265:14:freechips.rocketchip.system.DefaultConfig.fir@220375.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseeAck carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:266 assert (bundle.param === UInt(0), \"'D' channel ReleaseeAck carries invalid param\" + extra)\n"); // @[Monitor.scala 266:14:freechips.rocketchip.system.DefaultConfig.fir@220382.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 266:14:freechips.rocketchip.system.DefaultConfig.fir@220383.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:267 assert (!bundle.corrupt, \"'D' channel ReleaseAck is corrupt\" + extra)\n"); // @[Monitor.scala 267:14:freechips.rocketchip.system.DefaultConfig.fir@220390.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 267:14:freechips.rocketchip.system.DefaultConfig.fir@220391.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel ReleaseAck is denied (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:268 assert (!bundle.denied, \"'D' channel ReleaseAck is denied\" + extra)\n"); // @[Monitor.scala 268:14:freechips.rocketchip.system.DefaultConfig.fir@220398.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 268:14:freechips.rocketchip.system.DefaultConfig.fir@220399.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:272 assert (source_ok, \"'D' channel Grant carries invalid source ID\" + extra)\n"); // @[Monitor.scala 272:14:freechips.rocketchip.system.DefaultConfig.fir@220408.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 272:14:freechips.rocketchip.system.DefaultConfig.fir@220409.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid sink ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:273 assert (sink_ok, \"'D' channel Grant carries invalid sink ID\" + extra)\n"); // @[Monitor.scala 273:14:freechips.rocketchip.system.DefaultConfig.fir@220415.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_116) begin
          $fatal; // @[Monitor.scala 273:14:freechips.rocketchip.system.DefaultConfig.fir@220416.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_101 & _T_383) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant smaller than a beat (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:274 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel Grant smaller than a beat\" + extra)\n"); // @[Monitor.scala 274:14:freechips.rocketchip.system.DefaultConfig.fir@220423.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_101 & _T_383) begin
          $fatal; // @[Monitor.scala 274:14:freechips.rocketchip.system.DefaultConfig.fir@220424.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries invalid cap param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:275 assert (TLPermissions.isCap(bundle.param), \"'D' channel Grant carries invalid cap param\" + extra)\n"); // @[Monitor.scala 275:14:freechips.rocketchip.system.DefaultConfig.fir@220431.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 275:14:freechips.rocketchip.system.DefaultConfig.fir@220432.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant carries toN param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:276 assert (bundle.param =/= TLPermissions.toN, \"'D' channel Grant carries toN param\" + extra)\n"); // @[Monitor.scala 276:14:freechips.rocketchip.system.DefaultConfig.fir@220439.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 276:14:freechips.rocketchip.system.DefaultConfig.fir@220440.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:277 assert (!bundle.corrupt, \"'D' channel Grant is corrupt\" + extra)\n"); // @[Monitor.scala 277:14:freechips.rocketchip.system.DefaultConfig.fir@220447.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 277:14:freechips.rocketchip.system.DefaultConfig.fir@220448.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel Grant is denied (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:278 assert (deny_put_ok || !bundle.denied, \"'D' channel Grant is denied\" + extra)\n"); // @[Monitor.scala 278:14:freechips.rocketchip.system.DefaultConfig.fir@220456.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 278:14:freechips.rocketchip.system.DefaultConfig.fir@220457.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:282 assert (source_ok, \"'D' channel GrantData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 282:14:freechips.rocketchip.system.DefaultConfig.fir@220466.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 282:14:freechips.rocketchip.system.DefaultConfig.fir@220467.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_116) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid sink ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:283 assert (sink_ok, \"'D' channel GrantData carries invalid sink ID\" + extra)\n"); // @[Monitor.scala 283:14:freechips.rocketchip.system.DefaultConfig.fir@220473.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_116) begin
          $fatal; // @[Monitor.scala 283:14:freechips.rocketchip.system.DefaultConfig.fir@220474.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_105 & _T_383) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData smaller than a beat (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:284 assert (bundle.size >= UInt(log2Ceil(edge.manager.beatBytes)), \"'D' channel GrantData smaller than a beat\" + extra)\n"); // @[Monitor.scala 284:14:freechips.rocketchip.system.DefaultConfig.fir@220481.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_105 & _T_383) begin
          $fatal; // @[Monitor.scala 284:14:freechips.rocketchip.system.DefaultConfig.fir@220482.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries invalid cap param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:285 assert (TLPermissions.isCap(bundle.param), \"'D' channel GrantData carries invalid cap param\" + extra)\n"); // @[Monitor.scala 285:14:freechips.rocketchip.system.DefaultConfig.fir@220489.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 285:14:freechips.rocketchip.system.DefaultConfig.fir@220490.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData carries toN param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:286 assert (bundle.param =/= TLPermissions.toN, \"'D' channel GrantData carries toN param\" + extra)\n"); // @[Monitor.scala 286:14:freechips.rocketchip.system.DefaultConfig.fir@220497.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 286:14:freechips.rocketchip.system.DefaultConfig.fir@220498.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied but not corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:287 assert (!bundle.denied || bundle.corrupt, \"'D' channel GrantData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 287:14:freechips.rocketchip.system.DefaultConfig.fir@220506.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 287:14:freechips.rocketchip.system.DefaultConfig.fir@220507.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel GrantData is denied (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:288 assert (deny_get_ok || !bundle.denied, \"'D' channel GrantData is denied\" + extra)\n"); // @[Monitor.scala 288:14:freechips.rocketchip.system.DefaultConfig.fir@220515.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 288:14:freechips.rocketchip.system.DefaultConfig.fir@220516.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:292 assert (source_ok, \"'D' channel AccessAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 292:14:freechips.rocketchip.system.DefaultConfig.fir@220525.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 292:14:freechips.rocketchip.system.DefaultConfig.fir@220526.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:294 assert (bundle.param === UInt(0), \"'D' channel AccessAck carries invalid param\" + extra)\n"); // @[Monitor.scala 294:14:freechips.rocketchip.system.DefaultConfig.fir@220533.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 294:14:freechips.rocketchip.system.DefaultConfig.fir@220534.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:295 assert (!bundle.corrupt, \"'D' channel AccessAck is corrupt\" + extra)\n"); // @[Monitor.scala 295:14:freechips.rocketchip.system.DefaultConfig.fir@220541.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 295:14:freechips.rocketchip.system.DefaultConfig.fir@220542.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAck is denied (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:296 assert (deny_put_ok || !bundle.denied, \"'D' channel AccessAck is denied\" + extra)\n"); // @[Monitor.scala 296:14:freechips.rocketchip.system.DefaultConfig.fir@220550.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 296:14:freechips.rocketchip.system.DefaultConfig.fir@220551.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:300 assert (source_ok, \"'D' channel AccessAckData carries invalid source ID\" + extra)\n"); // @[Monitor.scala 300:14:freechips.rocketchip.system.DefaultConfig.fir@220560.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 300:14:freechips.rocketchip.system.DefaultConfig.fir@220561.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:302 assert (bundle.param === UInt(0), \"'D' channel AccessAckData carries invalid param\" + extra)\n"); // @[Monitor.scala 302:14:freechips.rocketchip.system.DefaultConfig.fir@220568.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 302:14:freechips.rocketchip.system.DefaultConfig.fir@220569.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied but not corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:303 assert (!bundle.denied || bundle.corrupt, \"'D' channel AccessAckData is denied but not corrupt\" + extra)\n"); // @[Monitor.scala 303:14:freechips.rocketchip.system.DefaultConfig.fir@220577.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 303:14:freechips.rocketchip.system.DefaultConfig.fir@220578.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel AccessAckData is denied (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:304 assert (deny_get_ok || !bundle.denied, \"'D' channel AccessAckData is denied\" + extra)\n"); // @[Monitor.scala 304:14:freechips.rocketchip.system.DefaultConfig.fir@220586.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 304:14:freechips.rocketchip.system.DefaultConfig.fir@220587.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:308 assert (source_ok, \"'D' channel HintAck carries invalid source ID\" + extra)\n"); // @[Monitor.scala 308:14:freechips.rocketchip.system.DefaultConfig.fir@220596.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 308:14:freechips.rocketchip.system.DefaultConfig.fir@220597.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck carries invalid param (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:310 assert (bundle.param === UInt(0), \"'D' channel HintAck carries invalid param\" + extra)\n"); // @[Monitor.scala 310:14:freechips.rocketchip.system.DefaultConfig.fir@220604.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 310:14:freechips.rocketchip.system.DefaultConfig.fir@220605.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is corrupt (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:311 assert (!bundle.corrupt, \"'D' channel HintAck is corrupt\" + extra)\n"); // @[Monitor.scala 311:14:freechips.rocketchip.system.DefaultConfig.fir@220612.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 311:14:freechips.rocketchip.system.DefaultConfig.fir@220613.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel HintAck is denied (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:312 assert (deny_put_ok || !bundle.denied, \"'D' channel HintAck is denied\" + extra)\n"); // @[Monitor.scala 312:14:freechips.rocketchip.system.DefaultConfig.fir@220621.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 312:14:freechips.rocketchip.system.DefaultConfig.fir@220622.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'B' channel valid and not TL-C (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:329 assert (!bundle.b.valid, \"'B' channel valid and not TL-C\" + extra)\n"); // @[Monitor.scala 329:14:freechips.rocketchip.system.DefaultConfig.fir@220631.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 329:14:freechips.rocketchip.system.DefaultConfig.fir@220632.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'C' channel valid and not TL-C (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:330 assert (!bundle.c.valid, \"'C' channel valid and not TL-C\" + extra)\n"); // @[Monitor.scala 330:14:freechips.rocketchip.system.DefaultConfig.fir@220639.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 330:14:freechips.rocketchip.system.DefaultConfig.fir@220640.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'E' channel valid and not TL-C (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:331 assert (!bundle.e.valid, \"'E' channel valid and not TL-C\" + extra)\n"); // @[Monitor.scala 331:14:freechips.rocketchip.system.DefaultConfig.fir@220647.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 331:14:freechips.rocketchip.system.DefaultConfig.fir@220648.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550 & _T_554) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel opcode changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:343 assert (a.bits.opcode === opcode, \"'A' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 343:14:freechips.rocketchip.system.DefaultConfig.fir@220687.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550 & _T_554) begin
          $fatal; // @[Monitor.scala 343:14:freechips.rocketchip.system.DefaultConfig.fir@220688.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550 & _T_558) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel param changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:344 assert (a.bits.param  === param,  \"'A' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 344:14:freechips.rocketchip.system.DefaultConfig.fir@220695.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550 & _T_558) begin
          $fatal; // @[Monitor.scala 344:14:freechips.rocketchip.system.DefaultConfig.fir@220696.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550 & _T_562) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel size changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:345 assert (a.bits.size   === size,   \"'A' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 345:14:freechips.rocketchip.system.DefaultConfig.fir@220703.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550 & _T_562) begin
          $fatal; // @[Monitor.scala 345:14:freechips.rocketchip.system.DefaultConfig.fir@220704.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550 & _T_566) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel source changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:346 assert (a.bits.source === source, \"'A' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 346:14:freechips.rocketchip.system.DefaultConfig.fir@220711.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550 & _T_566) begin
          $fatal; // @[Monitor.scala 346:14:freechips.rocketchip.system.DefaultConfig.fir@220712.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_550 & _T_570) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel address changed with multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:347 assert (a.bits.address=== address,\"'A' channel address changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 347:14:freechips.rocketchip.system.DefaultConfig.fir@220719.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_550 & _T_570) begin
          $fatal; // @[Monitor.scala 347:14:freechips.rocketchip.system.DefaultConfig.fir@220720.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_607 & _T_611) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel opcode changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:413 assert (d.bits.opcode === opcode, \"'D' channel opcode changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 413:14:freechips.rocketchip.system.DefaultConfig.fir@220769.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_607 & _T_611) begin
          $fatal; // @[Monitor.scala 413:14:freechips.rocketchip.system.DefaultConfig.fir@220770.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel param changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:414 assert (d.bits.param  === param,  \"'D' channel param changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 414:14:freechips.rocketchip.system.DefaultConfig.fir@220777.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 414:14:freechips.rocketchip.system.DefaultConfig.fir@220778.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_607 & _T_619) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel size changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:415 assert (d.bits.size   === size,   \"'D' channel size changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 415:14:freechips.rocketchip.system.DefaultConfig.fir@220785.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_607 & _T_619) begin
          $fatal; // @[Monitor.scala 415:14:freechips.rocketchip.system.DefaultConfig.fir@220786.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_607 & _T_623) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel source changed within multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:416 assert (d.bits.source === source, \"'D' channel source changed within multibeat operation\" + extra)\n"); // @[Monitor.scala 416:14:freechips.rocketchip.system.DefaultConfig.fir@220793.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_607 & _T_623) begin
          $fatal; // @[Monitor.scala 416:14:freechips.rocketchip.system.DefaultConfig.fir@220794.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel sink changed with multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:417 assert (d.bits.sink   === sink,   \"'D' channel sink changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 417:14:freechips.rocketchip.system.DefaultConfig.fir@220801.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 417:14:freechips.rocketchip.system.DefaultConfig.fir@220802.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel denied changed with multibeat operation (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:418 assert (d.bits.denied === denied, \"'D' channel denied changed with multibeat operation\" + extra)\n"); // @[Monitor.scala 418:14:freechips.rocketchip.system.DefaultConfig.fir@220809.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[Monitor.scala 418:14:freechips.rocketchip.system.DefaultConfig.fir@220810.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_682 & _T_690) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' channel re-used a source ID (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:448 assert(!inflight(bundle.a.bits.source), \"'A' channel re-used a source ID\" + extra)\n"); // @[Monitor.scala 448:13:freechips.rocketchip.system.DefaultConfig.fir@220887.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_682 & _T_690) begin
          $fatal; // @[Monitor.scala 448:13:freechips.rocketchip.system.DefaultConfig.fir@220888.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_698 & _T_705) begin
          $fwrite(32'h80000002,"Assertion failed: 'D' channel acknowledged for nothing inflight (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:455 assert((a_set | inflight)(bundle.d.bits.source), \"'D' channel acknowledged for nothing inflight\" + extra)\n"); // @[Monitor.scala 455:13:freechips.rocketchip.system.DefaultConfig.fir@220910.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_698 & _T_705) begin
          $fatal; // @[Monitor.scala 455:13:freechips.rocketchip.system.DefaultConfig.fir@220911.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_712) begin
          $fwrite(32'h80000002,"Assertion failed: 'A' and 'D' concurrent, despite minlatency 1 (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:459 assert(a_set =/= d_clr || !a_set.orR, s\"'A' and 'D' concurrent, despite minlatency ${edge.manager.minLatency}\" + extra)\n"); // @[Monitor.scala 459:13:freechips.rocketchip.system.DefaultConfig.fir@220922.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_712) begin
          $fatal; // @[Monitor.scala 459:13:freechips.rocketchip.system.DefaultConfig.fir@220923.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_726) begin
          $fwrite(32'h80000002,"Assertion failed: TileLink timeout expired (connected at MemoryBus.scala:80:46)\n    at Monitor.scala:467 assert (!inflight.orR || limit === UInt(0) || watchdog < limit, \"TileLink timeout expired\" + extra)\n"); // @[Monitor.scala 467:12:freechips.rocketchip.system.DefaultConfig.fir@220942.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_726) begin
          $fatal; // @[Monitor.scala 467:12:freechips.rocketchip.system.DefaultConfig.fir@220943.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
