module L2_meta_array(
  input  [10:0] RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input         RW0_wdata_0_valid,
  input         RW0_wdata_0_dirty,
  input  [15:0] RW0_wdata_0_tag,
  input         RW0_wdata_0_rr_state,
  input  [3:0]  RW0_wdata_0_dsid,
  input         RW0_wdata_1_valid,
  input         RW0_wdata_1_dirty,
  input  [15:0] RW0_wdata_1_tag,
  input         RW0_wdata_1_rr_state,
  input  [3:0]  RW0_wdata_1_dsid,
  input         RW0_wdata_2_valid,
  input         RW0_wdata_2_dirty,
  input  [15:0] RW0_wdata_2_tag,
  input         RW0_wdata_2_rr_state,
  input  [3:0]  RW0_wdata_2_dsid,
  input         RW0_wdata_3_valid,
  input         RW0_wdata_3_dirty,
  input  [15:0] RW0_wdata_3_tag,
  input         RW0_wdata_3_rr_state,
  input  [3:0]  RW0_wdata_3_dsid,
  input         RW0_wdata_4_valid,
  input         RW0_wdata_4_dirty,
  input  [15:0] RW0_wdata_4_tag,
  input         RW0_wdata_4_rr_state,
  input  [3:0]  RW0_wdata_4_dsid,
  input         RW0_wdata_5_valid,
  input         RW0_wdata_5_dirty,
  input  [15:0] RW0_wdata_5_tag,
  input         RW0_wdata_5_rr_state,
  input  [3:0]  RW0_wdata_5_dsid,
  input         RW0_wdata_6_valid,
  input         RW0_wdata_6_dirty,
  input  [15:0] RW0_wdata_6_tag,
  input         RW0_wdata_6_rr_state,
  input  [3:0]  RW0_wdata_6_dsid,
  input         RW0_wdata_7_valid,
  input         RW0_wdata_7_dirty,
  input  [15:0] RW0_wdata_7_tag,
  input         RW0_wdata_7_rr_state,
  input  [3:0]  RW0_wdata_7_dsid,
  input         RW0_wdata_8_valid,
  input         RW0_wdata_8_dirty,
  input  [15:0] RW0_wdata_8_tag,
  input         RW0_wdata_8_rr_state,
  input  [3:0]  RW0_wdata_8_dsid,
  input         RW0_wdata_9_valid,
  input         RW0_wdata_9_dirty,
  input  [15:0] RW0_wdata_9_tag,
  input         RW0_wdata_9_rr_state,
  input  [3:0]  RW0_wdata_9_dsid,
  input         RW0_wdata_10_valid,
  input         RW0_wdata_10_dirty,
  input  [15:0] RW0_wdata_10_tag,
  input         RW0_wdata_10_rr_state,
  input  [3:0]  RW0_wdata_10_dsid,
  input         RW0_wdata_11_valid,
  input         RW0_wdata_11_dirty,
  input  [15:0] RW0_wdata_11_tag,
  input         RW0_wdata_11_rr_state,
  input  [3:0]  RW0_wdata_11_dsid,
  input         RW0_wdata_12_valid,
  input         RW0_wdata_12_dirty,
  input  [15:0] RW0_wdata_12_tag,
  input         RW0_wdata_12_rr_state,
  input  [3:0]  RW0_wdata_12_dsid,
  input         RW0_wdata_13_valid,
  input         RW0_wdata_13_dirty,
  input  [15:0] RW0_wdata_13_tag,
  input         RW0_wdata_13_rr_state,
  input  [3:0]  RW0_wdata_13_dsid,
  input         RW0_wdata_14_valid,
  input         RW0_wdata_14_dirty,
  input  [15:0] RW0_wdata_14_tag,
  input         RW0_wdata_14_rr_state,
  input  [3:0]  RW0_wdata_14_dsid,
  input         RW0_wdata_15_valid,
  input         RW0_wdata_15_dirty,
  input  [15:0] RW0_wdata_15_tag,
  input         RW0_wdata_15_rr_state,
  input  [3:0]  RW0_wdata_15_dsid,
  output        RW0_rdata_0_valid,
  output        RW0_rdata_0_dirty,
  output [15:0] RW0_rdata_0_tag,
  output        RW0_rdata_0_rr_state,
  output [3:0]  RW0_rdata_0_dsid,
  output        RW0_rdata_1_valid,
  output        RW0_rdata_1_dirty,
  output [15:0] RW0_rdata_1_tag,
  output        RW0_rdata_1_rr_state,
  output [3:0]  RW0_rdata_1_dsid,
  output        RW0_rdata_2_valid,
  output        RW0_rdata_2_dirty,
  output [15:0] RW0_rdata_2_tag,
  output        RW0_rdata_2_rr_state,
  output [3:0]  RW0_rdata_2_dsid,
  output        RW0_rdata_3_valid,
  output        RW0_rdata_3_dirty,
  output [15:0] RW0_rdata_3_tag,
  output        RW0_rdata_3_rr_state,
  output [3:0]  RW0_rdata_3_dsid,
  output        RW0_rdata_4_valid,
  output        RW0_rdata_4_dirty,
  output [15:0] RW0_rdata_4_tag,
  output        RW0_rdata_4_rr_state,
  output [3:0]  RW0_rdata_4_dsid,
  output        RW0_rdata_5_valid,
  output        RW0_rdata_5_dirty,
  output [15:0] RW0_rdata_5_tag,
  output        RW0_rdata_5_rr_state,
  output [3:0]  RW0_rdata_5_dsid,
  output        RW0_rdata_6_valid,
  output        RW0_rdata_6_dirty,
  output [15:0] RW0_rdata_6_tag,
  output        RW0_rdata_6_rr_state,
  output [3:0]  RW0_rdata_6_dsid,
  output        RW0_rdata_7_valid,
  output        RW0_rdata_7_dirty,
  output [15:0] RW0_rdata_7_tag,
  output        RW0_rdata_7_rr_state,
  output [3:0]  RW0_rdata_7_dsid,
  output        RW0_rdata_8_valid,
  output        RW0_rdata_8_dirty,
  output [15:0] RW0_rdata_8_tag,
  output        RW0_rdata_8_rr_state,
  output [3:0]  RW0_rdata_8_dsid,
  output        RW0_rdata_9_valid,
  output        RW0_rdata_9_dirty,
  output [15:0] RW0_rdata_9_tag,
  output        RW0_rdata_9_rr_state,
  output [3:0]  RW0_rdata_9_dsid,
  output        RW0_rdata_10_valid,
  output        RW0_rdata_10_dirty,
  output [15:0] RW0_rdata_10_tag,
  output        RW0_rdata_10_rr_state,
  output [3:0]  RW0_rdata_10_dsid,
  output        RW0_rdata_11_valid,
  output        RW0_rdata_11_dirty,
  output [15:0] RW0_rdata_11_tag,
  output        RW0_rdata_11_rr_state,
  output [3:0]  RW0_rdata_11_dsid,
  output        RW0_rdata_12_valid,
  output        RW0_rdata_12_dirty,
  output [15:0] RW0_rdata_12_tag,
  output        RW0_rdata_12_rr_state,
  output [3:0]  RW0_rdata_12_dsid,
  output        RW0_rdata_13_valid,
  output        RW0_rdata_13_dirty,
  output [15:0] RW0_rdata_13_tag,
  output        RW0_rdata_13_rr_state,
  output [3:0]  RW0_rdata_13_dsid,
  output        RW0_rdata_14_valid,
  output        RW0_rdata_14_dirty,
  output [15:0] RW0_rdata_14_tag,
  output        RW0_rdata_14_rr_state,
  output [3:0]  RW0_rdata_14_dsid,
  output        RW0_rdata_15_valid,
  output        RW0_rdata_15_dirty,
  output [15:0] RW0_rdata_15_tag,
  output        RW0_rdata_15_rr_state,
  output [3:0]  RW0_rdata_15_dsid
);
  wire [10:0] L2_meta_array_ext_RW0_addr;
  wire  L2_meta_array_ext_RW0_en;
  wire  L2_meta_array_ext_RW0_clk;
  wire  L2_meta_array_ext_RW0_wmode;
  wire [367:0] L2_meta_array_ext_RW0_wdata;
  wire [367:0] L2_meta_array_ext_RW0_rdata;
  wire [3:0] _GEN_0;
  wire  _GEN_1;
  wire [15:0] _GEN_2;
  wire  _GEN_3;
  wire  _GEN_4;
  wire [3:0] _GEN_5;
  wire  _GEN_6;
  wire [15:0] _GEN_7;
  wire  _GEN_8;
  wire  _GEN_9;
  wire [3:0] _GEN_10;
  wire  _GEN_11;
  wire [15:0] _GEN_12;
  wire  _GEN_13;
  wire  _GEN_14;
  wire [3:0] _GEN_15;
  wire  _GEN_16;
  wire [15:0] _GEN_17;
  wire  _GEN_18;
  wire  _GEN_19;
  wire [3:0] _GEN_20;
  wire  _GEN_21;
  wire [15:0] _GEN_22;
  wire  _GEN_23;
  wire  _GEN_24;
  wire [3:0] _GEN_25;
  wire  _GEN_26;
  wire [15:0] _GEN_27;
  wire  _GEN_28;
  wire  _GEN_29;
  wire [3:0] _GEN_30;
  wire  _GEN_31;
  wire [15:0] _GEN_32;
  wire  _GEN_33;
  wire  _GEN_34;
  wire [3:0] _GEN_35;
  wire  _GEN_36;
  wire [15:0] _GEN_37;
  wire  _GEN_38;
  wire  _GEN_39;
  wire [3:0] _GEN_40;
  wire  _GEN_41;
  wire [15:0] _GEN_42;
  wire  _GEN_43;
  wire  _GEN_44;
  wire [3:0] _GEN_45;
  wire  _GEN_46;
  wire [15:0] _GEN_47;
  wire  _GEN_48;
  wire  _GEN_49;
  wire [3:0] _GEN_50;
  wire  _GEN_51;
  wire [15:0] _GEN_52;
  wire  _GEN_53;
  wire  _GEN_54;
  wire [3:0] _GEN_55;
  wire  _GEN_56;
  wire [15:0] _GEN_57;
  wire  _GEN_58;
  wire  _GEN_59;
  wire [3:0] _GEN_60;
  wire  _GEN_61;
  wire [15:0] _GEN_62;
  wire  _GEN_63;
  wire  _GEN_64;
  wire [3:0] _GEN_65;
  wire  _GEN_66;
  wire [15:0] _GEN_67;
  wire  _GEN_68;
  wire  _GEN_69;
  wire [3:0] _GEN_70;
  wire  _GEN_71;
  wire [15:0] _GEN_72;
  wire  _GEN_73;
  wire  _GEN_74;
  wire [3:0] _GEN_75;
  wire  _GEN_76;
  wire [15:0] _GEN_77;
  wire  _GEN_78;
  wire  _GEN_79;
  wire  _GEN_80;
  wire  _GEN_81;
  wire  _GEN_82;
  wire [3:0] _GEN_83;
  wire [15:0] _GEN_84;
  wire [4:0] _GEN_85;
  wire [1:0] _GEN_86;
  wire [20:0] _GEN_87;
  wire  _GEN_88;
  wire  _GEN_89;
  wire  _GEN_90;
  wire [3:0] _GEN_91;
  wire [15:0] _GEN_92;
  wire [4:0] _GEN_93;
  wire [1:0] _GEN_94;
  wire [20:0] _GEN_95;
  wire [22:0] _GEN_96;
  wire [22:0] _GEN_97;
  wire  _GEN_98;
  wire  _GEN_99;
  wire  _GEN_100;
  wire [3:0] _GEN_101;
  wire [15:0] _GEN_102;
  wire [4:0] _GEN_103;
  wire [1:0] _GEN_104;
  wire [20:0] _GEN_105;
  wire  _GEN_106;
  wire  _GEN_107;
  wire  _GEN_108;
  wire [3:0] _GEN_109;
  wire [15:0] _GEN_110;
  wire [4:0] _GEN_111;
  wire [1:0] _GEN_112;
  wire [20:0] _GEN_113;
  wire [22:0] _GEN_114;
  wire [22:0] _GEN_115;
  wire [45:0] _GEN_116;
  wire [45:0] _GEN_117;
  wire  _GEN_118;
  wire  _GEN_119;
  wire  _GEN_120;
  wire [3:0] _GEN_121;
  wire [15:0] _GEN_122;
  wire [4:0] _GEN_123;
  wire [1:0] _GEN_124;
  wire [20:0] _GEN_125;
  wire  _GEN_126;
  wire  _GEN_127;
  wire  _GEN_128;
  wire [3:0] _GEN_129;
  wire [15:0] _GEN_130;
  wire [4:0] _GEN_131;
  wire [1:0] _GEN_132;
  wire [20:0] _GEN_133;
  wire [22:0] _GEN_134;
  wire [22:0] _GEN_135;
  wire  _GEN_136;
  wire  _GEN_137;
  wire  _GEN_138;
  wire [3:0] _GEN_139;
  wire [15:0] _GEN_140;
  wire [4:0] _GEN_141;
  wire [1:0] _GEN_142;
  wire [20:0] _GEN_143;
  wire  _GEN_144;
  wire  _GEN_145;
  wire  _GEN_146;
  wire [3:0] _GEN_147;
  wire [15:0] _GEN_148;
  wire [4:0] _GEN_149;
  wire [1:0] _GEN_150;
  wire [20:0] _GEN_151;
  wire [22:0] _GEN_152;
  wire [22:0] _GEN_153;
  wire [45:0] _GEN_154;
  wire [45:0] _GEN_155;
  wire [91:0] _GEN_156;
  wire [91:0] _GEN_157;
  wire  _GEN_158;
  wire  _GEN_159;
  wire  _GEN_160;
  wire [3:0] _GEN_161;
  wire [15:0] _GEN_162;
  wire [4:0] _GEN_163;
  wire [1:0] _GEN_164;
  wire [20:0] _GEN_165;
  wire  _GEN_166;
  wire  _GEN_167;
  wire  _GEN_168;
  wire [3:0] _GEN_169;
  wire [15:0] _GEN_170;
  wire [4:0] _GEN_171;
  wire [1:0] _GEN_172;
  wire [20:0] _GEN_173;
  wire [22:0] _GEN_174;
  wire [22:0] _GEN_175;
  wire  _GEN_176;
  wire  _GEN_177;
  wire  _GEN_178;
  wire [3:0] _GEN_179;
  wire [15:0] _GEN_180;
  wire [4:0] _GEN_181;
  wire [1:0] _GEN_182;
  wire [20:0] _GEN_183;
  wire  _GEN_184;
  wire  _GEN_185;
  wire  _GEN_186;
  wire [3:0] _GEN_187;
  wire [15:0] _GEN_188;
  wire [4:0] _GEN_189;
  wire [1:0] _GEN_190;
  wire [20:0] _GEN_191;
  wire [22:0] _GEN_192;
  wire [22:0] _GEN_193;
  wire [45:0] _GEN_194;
  wire [45:0] _GEN_195;
  wire  _GEN_196;
  wire  _GEN_197;
  wire  _GEN_198;
  wire [3:0] _GEN_199;
  wire [15:0] _GEN_200;
  wire [4:0] _GEN_201;
  wire [1:0] _GEN_202;
  wire [20:0] _GEN_203;
  wire  _GEN_204;
  wire  _GEN_205;
  wire  _GEN_206;
  wire [3:0] _GEN_207;
  wire [15:0] _GEN_208;
  wire [4:0] _GEN_209;
  wire [1:0] _GEN_210;
  wire [20:0] _GEN_211;
  wire [22:0] _GEN_212;
  wire [22:0] _GEN_213;
  wire  _GEN_214;
  wire  _GEN_215;
  wire  _GEN_216;
  wire [3:0] _GEN_217;
  wire [15:0] _GEN_218;
  wire [4:0] _GEN_219;
  wire [1:0] _GEN_220;
  wire [20:0] _GEN_221;
  wire  _GEN_222;
  wire  _GEN_223;
  wire  _GEN_224;
  wire [3:0] _GEN_225;
  wire [15:0] _GEN_226;
  wire [4:0] _GEN_227;
  wire [1:0] _GEN_228;
  wire [20:0] _GEN_229;
  wire [22:0] _GEN_230;
  wire [22:0] _GEN_231;
  wire [45:0] _GEN_232;
  wire [45:0] _GEN_233;
  wire [91:0] _GEN_234;
  wire [91:0] _GEN_235;
  wire [183:0] _GEN_236;
  wire [183:0] _GEN_237;
  L2_meta_array_ext L2_meta_array_ext (
    .RW0_addr(L2_meta_array_ext_RW0_addr),
    .RW0_en(L2_meta_array_ext_RW0_en),
    .RW0_clk(L2_meta_array_ext_RW0_clk),
    .RW0_wmode(L2_meta_array_ext_RW0_wmode),
    .RW0_wdata(L2_meta_array_ext_RW0_wdata),
    .RW0_rdata(L2_meta_array_ext_RW0_rdata)
  );
  assign L2_meta_array_ext_RW0_clk = RW0_clk;
  assign L2_meta_array_ext_RW0_en = RW0_en;
  assign L2_meta_array_ext_RW0_addr = RW0_addr;
  assign _GEN_0 = L2_meta_array_ext_RW0_rdata[3:0];
  assign RW0_rdata_0_dsid = $unsigned(_GEN_0);
  assign _GEN_1 = L2_meta_array_ext_RW0_rdata[4];
  assign RW0_rdata_0_rr_state = $unsigned(_GEN_1);
  assign _GEN_2 = L2_meta_array_ext_RW0_rdata[20:5];
  assign RW0_rdata_0_tag = $unsigned(_GEN_2);
  assign _GEN_3 = L2_meta_array_ext_RW0_rdata[21];
  assign RW0_rdata_0_dirty = $unsigned(_GEN_3);
  assign _GEN_4 = L2_meta_array_ext_RW0_rdata[22];
  assign RW0_rdata_0_valid = $unsigned(_GEN_4);
  assign _GEN_5 = L2_meta_array_ext_RW0_rdata[26:23];
  assign RW0_rdata_1_dsid = $unsigned(_GEN_5);
  assign _GEN_6 = L2_meta_array_ext_RW0_rdata[27];
  assign RW0_rdata_1_rr_state = $unsigned(_GEN_6);
  assign _GEN_7 = L2_meta_array_ext_RW0_rdata[43:28];
  assign RW0_rdata_1_tag = $unsigned(_GEN_7);
  assign _GEN_8 = L2_meta_array_ext_RW0_rdata[44];
  assign RW0_rdata_1_dirty = $unsigned(_GEN_8);
  assign _GEN_9 = L2_meta_array_ext_RW0_rdata[45];
  assign RW0_rdata_1_valid = $unsigned(_GEN_9);
  assign _GEN_10 = L2_meta_array_ext_RW0_rdata[49:46];
  assign RW0_rdata_2_dsid = $unsigned(_GEN_10);
  assign _GEN_11 = L2_meta_array_ext_RW0_rdata[50];
  assign RW0_rdata_2_rr_state = $unsigned(_GEN_11);
  assign _GEN_12 = L2_meta_array_ext_RW0_rdata[66:51];
  assign RW0_rdata_2_tag = $unsigned(_GEN_12);
  assign _GEN_13 = L2_meta_array_ext_RW0_rdata[67];
  assign RW0_rdata_2_dirty = $unsigned(_GEN_13);
  assign _GEN_14 = L2_meta_array_ext_RW0_rdata[68];
  assign RW0_rdata_2_valid = $unsigned(_GEN_14);
  assign _GEN_15 = L2_meta_array_ext_RW0_rdata[72:69];
  assign RW0_rdata_3_dsid = $unsigned(_GEN_15);
  assign _GEN_16 = L2_meta_array_ext_RW0_rdata[73];
  assign RW0_rdata_3_rr_state = $unsigned(_GEN_16);
  assign _GEN_17 = L2_meta_array_ext_RW0_rdata[89:74];
  assign RW0_rdata_3_tag = $unsigned(_GEN_17);
  assign _GEN_18 = L2_meta_array_ext_RW0_rdata[90];
  assign RW0_rdata_3_dirty = $unsigned(_GEN_18);
  assign _GEN_19 = L2_meta_array_ext_RW0_rdata[91];
  assign RW0_rdata_3_valid = $unsigned(_GEN_19);
  assign _GEN_20 = L2_meta_array_ext_RW0_rdata[95:92];
  assign RW0_rdata_4_dsid = $unsigned(_GEN_20);
  assign _GEN_21 = L2_meta_array_ext_RW0_rdata[96];
  assign RW0_rdata_4_rr_state = $unsigned(_GEN_21);
  assign _GEN_22 = L2_meta_array_ext_RW0_rdata[112:97];
  assign RW0_rdata_4_tag = $unsigned(_GEN_22);
  assign _GEN_23 = L2_meta_array_ext_RW0_rdata[113];
  assign RW0_rdata_4_dirty = $unsigned(_GEN_23);
  assign _GEN_24 = L2_meta_array_ext_RW0_rdata[114];
  assign RW0_rdata_4_valid = $unsigned(_GEN_24);
  assign _GEN_25 = L2_meta_array_ext_RW0_rdata[118:115];
  assign RW0_rdata_5_dsid = $unsigned(_GEN_25);
  assign _GEN_26 = L2_meta_array_ext_RW0_rdata[119];
  assign RW0_rdata_5_rr_state = $unsigned(_GEN_26);
  assign _GEN_27 = L2_meta_array_ext_RW0_rdata[135:120];
  assign RW0_rdata_5_tag = $unsigned(_GEN_27);
  assign _GEN_28 = L2_meta_array_ext_RW0_rdata[136];
  assign RW0_rdata_5_dirty = $unsigned(_GEN_28);
  assign _GEN_29 = L2_meta_array_ext_RW0_rdata[137];
  assign RW0_rdata_5_valid = $unsigned(_GEN_29);
  assign _GEN_30 = L2_meta_array_ext_RW0_rdata[141:138];
  assign RW0_rdata_6_dsid = $unsigned(_GEN_30);
  assign _GEN_31 = L2_meta_array_ext_RW0_rdata[142];
  assign RW0_rdata_6_rr_state = $unsigned(_GEN_31);
  assign _GEN_32 = L2_meta_array_ext_RW0_rdata[158:143];
  assign RW0_rdata_6_tag = $unsigned(_GEN_32);
  assign _GEN_33 = L2_meta_array_ext_RW0_rdata[159];
  assign RW0_rdata_6_dirty = $unsigned(_GEN_33);
  assign _GEN_34 = L2_meta_array_ext_RW0_rdata[160];
  assign RW0_rdata_6_valid = $unsigned(_GEN_34);
  assign _GEN_35 = L2_meta_array_ext_RW0_rdata[164:161];
  assign RW0_rdata_7_dsid = $unsigned(_GEN_35);
  assign _GEN_36 = L2_meta_array_ext_RW0_rdata[165];
  assign RW0_rdata_7_rr_state = $unsigned(_GEN_36);
  assign _GEN_37 = L2_meta_array_ext_RW0_rdata[181:166];
  assign RW0_rdata_7_tag = $unsigned(_GEN_37);
  assign _GEN_38 = L2_meta_array_ext_RW0_rdata[182];
  assign RW0_rdata_7_dirty = $unsigned(_GEN_38);
  assign _GEN_39 = L2_meta_array_ext_RW0_rdata[183];
  assign RW0_rdata_7_valid = $unsigned(_GEN_39);
  assign _GEN_40 = L2_meta_array_ext_RW0_rdata[187:184];
  assign RW0_rdata_8_dsid = $unsigned(_GEN_40);
  assign _GEN_41 = L2_meta_array_ext_RW0_rdata[188];
  assign RW0_rdata_8_rr_state = $unsigned(_GEN_41);
  assign _GEN_42 = L2_meta_array_ext_RW0_rdata[204:189];
  assign RW0_rdata_8_tag = $unsigned(_GEN_42);
  assign _GEN_43 = L2_meta_array_ext_RW0_rdata[205];
  assign RW0_rdata_8_dirty = $unsigned(_GEN_43);
  assign _GEN_44 = L2_meta_array_ext_RW0_rdata[206];
  assign RW0_rdata_8_valid = $unsigned(_GEN_44);
  assign _GEN_45 = L2_meta_array_ext_RW0_rdata[210:207];
  assign RW0_rdata_9_dsid = $unsigned(_GEN_45);
  assign _GEN_46 = L2_meta_array_ext_RW0_rdata[211];
  assign RW0_rdata_9_rr_state = $unsigned(_GEN_46);
  assign _GEN_47 = L2_meta_array_ext_RW0_rdata[227:212];
  assign RW0_rdata_9_tag = $unsigned(_GEN_47);
  assign _GEN_48 = L2_meta_array_ext_RW0_rdata[228];
  assign RW0_rdata_9_dirty = $unsigned(_GEN_48);
  assign _GEN_49 = L2_meta_array_ext_RW0_rdata[229];
  assign RW0_rdata_9_valid = $unsigned(_GEN_49);
  assign _GEN_50 = L2_meta_array_ext_RW0_rdata[233:230];
  assign RW0_rdata_10_dsid = $unsigned(_GEN_50);
  assign _GEN_51 = L2_meta_array_ext_RW0_rdata[234];
  assign RW0_rdata_10_rr_state = $unsigned(_GEN_51);
  assign _GEN_52 = L2_meta_array_ext_RW0_rdata[250:235];
  assign RW0_rdata_10_tag = $unsigned(_GEN_52);
  assign _GEN_53 = L2_meta_array_ext_RW0_rdata[251];
  assign RW0_rdata_10_dirty = $unsigned(_GEN_53);
  assign _GEN_54 = L2_meta_array_ext_RW0_rdata[252];
  assign RW0_rdata_10_valid = $unsigned(_GEN_54);
  assign _GEN_55 = L2_meta_array_ext_RW0_rdata[256:253];
  assign RW0_rdata_11_dsid = $unsigned(_GEN_55);
  assign _GEN_56 = L2_meta_array_ext_RW0_rdata[257];
  assign RW0_rdata_11_rr_state = $unsigned(_GEN_56);
  assign _GEN_57 = L2_meta_array_ext_RW0_rdata[273:258];
  assign RW0_rdata_11_tag = $unsigned(_GEN_57);
  assign _GEN_58 = L2_meta_array_ext_RW0_rdata[274];
  assign RW0_rdata_11_dirty = $unsigned(_GEN_58);
  assign _GEN_59 = L2_meta_array_ext_RW0_rdata[275];
  assign RW0_rdata_11_valid = $unsigned(_GEN_59);
  assign _GEN_60 = L2_meta_array_ext_RW0_rdata[279:276];
  assign RW0_rdata_12_dsid = $unsigned(_GEN_60);
  assign _GEN_61 = L2_meta_array_ext_RW0_rdata[280];
  assign RW0_rdata_12_rr_state = $unsigned(_GEN_61);
  assign _GEN_62 = L2_meta_array_ext_RW0_rdata[296:281];
  assign RW0_rdata_12_tag = $unsigned(_GEN_62);
  assign _GEN_63 = L2_meta_array_ext_RW0_rdata[297];
  assign RW0_rdata_12_dirty = $unsigned(_GEN_63);
  assign _GEN_64 = L2_meta_array_ext_RW0_rdata[298];
  assign RW0_rdata_12_valid = $unsigned(_GEN_64);
  assign _GEN_65 = L2_meta_array_ext_RW0_rdata[302:299];
  assign RW0_rdata_13_dsid = $unsigned(_GEN_65);
  assign _GEN_66 = L2_meta_array_ext_RW0_rdata[303];
  assign RW0_rdata_13_rr_state = $unsigned(_GEN_66);
  assign _GEN_67 = L2_meta_array_ext_RW0_rdata[319:304];
  assign RW0_rdata_13_tag = $unsigned(_GEN_67);
  assign _GEN_68 = L2_meta_array_ext_RW0_rdata[320];
  assign RW0_rdata_13_dirty = $unsigned(_GEN_68);
  assign _GEN_69 = L2_meta_array_ext_RW0_rdata[321];
  assign RW0_rdata_13_valid = $unsigned(_GEN_69);
  assign _GEN_70 = L2_meta_array_ext_RW0_rdata[325:322];
  assign RW0_rdata_14_dsid = $unsigned(_GEN_70);
  assign _GEN_71 = L2_meta_array_ext_RW0_rdata[326];
  assign RW0_rdata_14_rr_state = $unsigned(_GEN_71);
  assign _GEN_72 = L2_meta_array_ext_RW0_rdata[342:327];
  assign RW0_rdata_14_tag = $unsigned(_GEN_72);
  assign _GEN_73 = L2_meta_array_ext_RW0_rdata[343];
  assign RW0_rdata_14_dirty = $unsigned(_GEN_73);
  assign _GEN_74 = L2_meta_array_ext_RW0_rdata[344];
  assign RW0_rdata_14_valid = $unsigned(_GEN_74);
  assign _GEN_75 = L2_meta_array_ext_RW0_rdata[348:345];
  assign RW0_rdata_15_dsid = $unsigned(_GEN_75);
  assign _GEN_76 = L2_meta_array_ext_RW0_rdata[349];
  assign RW0_rdata_15_rr_state = $unsigned(_GEN_76);
  assign _GEN_77 = L2_meta_array_ext_RW0_rdata[365:350];
  assign RW0_rdata_15_tag = $unsigned(_GEN_77);
  assign _GEN_78 = L2_meta_array_ext_RW0_rdata[366];
  assign RW0_rdata_15_dirty = $unsigned(_GEN_78);
  assign _GEN_79 = L2_meta_array_ext_RW0_rdata[367];
  assign RW0_rdata_15_valid = $unsigned(_GEN_79);
  assign L2_meta_array_ext_RW0_wmode = RW0_wmode;
  assign _GEN_80 = $unsigned(RW0_wdata_15_valid);
  assign _GEN_81 = $unsigned(RW0_wdata_15_dirty);
  assign _GEN_82 = $unsigned(RW0_wdata_15_rr_state);
  assign _GEN_83 = $unsigned(RW0_wdata_15_dsid);
  assign _GEN_84 = $unsigned(RW0_wdata_15_tag);
  assign _GEN_85 = {_GEN_82,_GEN_83};
  assign _GEN_86 = {_GEN_80,_GEN_81};
  assign _GEN_87 = {_GEN_84,_GEN_85};
  assign _GEN_88 = $unsigned(RW0_wdata_14_valid);
  assign _GEN_89 = $unsigned(RW0_wdata_14_dirty);
  assign _GEN_90 = $unsigned(RW0_wdata_14_rr_state);
  assign _GEN_91 = $unsigned(RW0_wdata_14_dsid);
  assign _GEN_92 = $unsigned(RW0_wdata_14_tag);
  assign _GEN_93 = {_GEN_90,_GEN_91};
  assign _GEN_94 = {_GEN_88,_GEN_89};
  assign _GEN_95 = {_GEN_92,_GEN_93};
  assign _GEN_96 = {_GEN_86,_GEN_87};
  assign _GEN_97 = {_GEN_94,_GEN_95};
  assign _GEN_98 = $unsigned(RW0_wdata_13_valid);
  assign _GEN_99 = $unsigned(RW0_wdata_13_dirty);
  assign _GEN_100 = $unsigned(RW0_wdata_13_rr_state);
  assign _GEN_101 = $unsigned(RW0_wdata_13_dsid);
  assign _GEN_102 = $unsigned(RW0_wdata_13_tag);
  assign _GEN_103 = {_GEN_100,_GEN_101};
  assign _GEN_104 = {_GEN_98,_GEN_99};
  assign _GEN_105 = {_GEN_102,_GEN_103};
  assign _GEN_106 = $unsigned(RW0_wdata_12_valid);
  assign _GEN_107 = $unsigned(RW0_wdata_12_dirty);
  assign _GEN_108 = $unsigned(RW0_wdata_12_rr_state);
  assign _GEN_109 = $unsigned(RW0_wdata_12_dsid);
  assign _GEN_110 = $unsigned(RW0_wdata_12_tag);
  assign _GEN_111 = {_GEN_108,_GEN_109};
  assign _GEN_112 = {_GEN_106,_GEN_107};
  assign _GEN_113 = {_GEN_110,_GEN_111};
  assign _GEN_114 = {_GEN_104,_GEN_105};
  assign _GEN_115 = {_GEN_112,_GEN_113};
  assign _GEN_116 = {_GEN_96,_GEN_97};
  assign _GEN_117 = {_GEN_114,_GEN_115};
  assign _GEN_118 = $unsigned(RW0_wdata_11_valid);
  assign _GEN_119 = $unsigned(RW0_wdata_11_dirty);
  assign _GEN_120 = $unsigned(RW0_wdata_11_rr_state);
  assign _GEN_121 = $unsigned(RW0_wdata_11_dsid);
  assign _GEN_122 = $unsigned(RW0_wdata_11_tag);
  assign _GEN_123 = {_GEN_120,_GEN_121};
  assign _GEN_124 = {_GEN_118,_GEN_119};
  assign _GEN_125 = {_GEN_122,_GEN_123};
  assign _GEN_126 = $unsigned(RW0_wdata_10_valid);
  assign _GEN_127 = $unsigned(RW0_wdata_10_dirty);
  assign _GEN_128 = $unsigned(RW0_wdata_10_rr_state);
  assign _GEN_129 = $unsigned(RW0_wdata_10_dsid);
  assign _GEN_130 = $unsigned(RW0_wdata_10_tag);
  assign _GEN_131 = {_GEN_128,_GEN_129};
  assign _GEN_132 = {_GEN_126,_GEN_127};
  assign _GEN_133 = {_GEN_130,_GEN_131};
  assign _GEN_134 = {_GEN_124,_GEN_125};
  assign _GEN_135 = {_GEN_132,_GEN_133};
  assign _GEN_136 = $unsigned(RW0_wdata_9_valid);
  assign _GEN_137 = $unsigned(RW0_wdata_9_dirty);
  assign _GEN_138 = $unsigned(RW0_wdata_9_rr_state);
  assign _GEN_139 = $unsigned(RW0_wdata_9_dsid);
  assign _GEN_140 = $unsigned(RW0_wdata_9_tag);
  assign _GEN_141 = {_GEN_138,_GEN_139};
  assign _GEN_142 = {_GEN_136,_GEN_137};
  assign _GEN_143 = {_GEN_140,_GEN_141};
  assign _GEN_144 = $unsigned(RW0_wdata_8_valid);
  assign _GEN_145 = $unsigned(RW0_wdata_8_dirty);
  assign _GEN_146 = $unsigned(RW0_wdata_8_rr_state);
  assign _GEN_147 = $unsigned(RW0_wdata_8_dsid);
  assign _GEN_148 = $unsigned(RW0_wdata_8_tag);
  assign _GEN_149 = {_GEN_146,_GEN_147};
  assign _GEN_150 = {_GEN_144,_GEN_145};
  assign _GEN_151 = {_GEN_148,_GEN_149};
  assign _GEN_152 = {_GEN_142,_GEN_143};
  assign _GEN_153 = {_GEN_150,_GEN_151};
  assign _GEN_154 = {_GEN_134,_GEN_135};
  assign _GEN_155 = {_GEN_152,_GEN_153};
  assign _GEN_156 = {_GEN_116,_GEN_117};
  assign _GEN_157 = {_GEN_154,_GEN_155};
  assign _GEN_158 = $unsigned(RW0_wdata_7_valid);
  assign _GEN_159 = $unsigned(RW0_wdata_7_dirty);
  assign _GEN_160 = $unsigned(RW0_wdata_7_rr_state);
  assign _GEN_161 = $unsigned(RW0_wdata_7_dsid);
  assign _GEN_162 = $unsigned(RW0_wdata_7_tag);
  assign _GEN_163 = {_GEN_160,_GEN_161};
  assign _GEN_164 = {_GEN_158,_GEN_159};
  assign _GEN_165 = {_GEN_162,_GEN_163};
  assign _GEN_166 = $unsigned(RW0_wdata_6_valid);
  assign _GEN_167 = $unsigned(RW0_wdata_6_dirty);
  assign _GEN_168 = $unsigned(RW0_wdata_6_rr_state);
  assign _GEN_169 = $unsigned(RW0_wdata_6_dsid);
  assign _GEN_170 = $unsigned(RW0_wdata_6_tag);
  assign _GEN_171 = {_GEN_168,_GEN_169};
  assign _GEN_172 = {_GEN_166,_GEN_167};
  assign _GEN_173 = {_GEN_170,_GEN_171};
  assign _GEN_174 = {_GEN_164,_GEN_165};
  assign _GEN_175 = {_GEN_172,_GEN_173};
  assign _GEN_176 = $unsigned(RW0_wdata_5_valid);
  assign _GEN_177 = $unsigned(RW0_wdata_5_dirty);
  assign _GEN_178 = $unsigned(RW0_wdata_5_rr_state);
  assign _GEN_179 = $unsigned(RW0_wdata_5_dsid);
  assign _GEN_180 = $unsigned(RW0_wdata_5_tag);
  assign _GEN_181 = {_GEN_178,_GEN_179};
  assign _GEN_182 = {_GEN_176,_GEN_177};
  assign _GEN_183 = {_GEN_180,_GEN_181};
  assign _GEN_184 = $unsigned(RW0_wdata_4_valid);
  assign _GEN_185 = $unsigned(RW0_wdata_4_dirty);
  assign _GEN_186 = $unsigned(RW0_wdata_4_rr_state);
  assign _GEN_187 = $unsigned(RW0_wdata_4_dsid);
  assign _GEN_188 = $unsigned(RW0_wdata_4_tag);
  assign _GEN_189 = {_GEN_186,_GEN_187};
  assign _GEN_190 = {_GEN_184,_GEN_185};
  assign _GEN_191 = {_GEN_188,_GEN_189};
  assign _GEN_192 = {_GEN_182,_GEN_183};
  assign _GEN_193 = {_GEN_190,_GEN_191};
  assign _GEN_194 = {_GEN_174,_GEN_175};
  assign _GEN_195 = {_GEN_192,_GEN_193};
  assign _GEN_196 = $unsigned(RW0_wdata_3_valid);
  assign _GEN_197 = $unsigned(RW0_wdata_3_dirty);
  assign _GEN_198 = $unsigned(RW0_wdata_3_rr_state);
  assign _GEN_199 = $unsigned(RW0_wdata_3_dsid);
  assign _GEN_200 = $unsigned(RW0_wdata_3_tag);
  assign _GEN_201 = {_GEN_198,_GEN_199};
  assign _GEN_202 = {_GEN_196,_GEN_197};
  assign _GEN_203 = {_GEN_200,_GEN_201};
  assign _GEN_204 = $unsigned(RW0_wdata_2_valid);
  assign _GEN_205 = $unsigned(RW0_wdata_2_dirty);
  assign _GEN_206 = $unsigned(RW0_wdata_2_rr_state);
  assign _GEN_207 = $unsigned(RW0_wdata_2_dsid);
  assign _GEN_208 = $unsigned(RW0_wdata_2_tag);
  assign _GEN_209 = {_GEN_206,_GEN_207};
  assign _GEN_210 = {_GEN_204,_GEN_205};
  assign _GEN_211 = {_GEN_208,_GEN_209};
  assign _GEN_212 = {_GEN_202,_GEN_203};
  assign _GEN_213 = {_GEN_210,_GEN_211};
  assign _GEN_214 = $unsigned(RW0_wdata_1_valid);
  assign _GEN_215 = $unsigned(RW0_wdata_1_dirty);
  assign _GEN_216 = $unsigned(RW0_wdata_1_rr_state);
  assign _GEN_217 = $unsigned(RW0_wdata_1_dsid);
  assign _GEN_218 = $unsigned(RW0_wdata_1_tag);
  assign _GEN_219 = {_GEN_216,_GEN_217};
  assign _GEN_220 = {_GEN_214,_GEN_215};
  assign _GEN_221 = {_GEN_218,_GEN_219};
  assign _GEN_222 = $unsigned(RW0_wdata_0_valid);
  assign _GEN_223 = $unsigned(RW0_wdata_0_dirty);
  assign _GEN_224 = $unsigned(RW0_wdata_0_rr_state);
  assign _GEN_225 = $unsigned(RW0_wdata_0_dsid);
  assign _GEN_226 = $unsigned(RW0_wdata_0_tag);
  assign _GEN_227 = {_GEN_224,_GEN_225};
  assign _GEN_228 = {_GEN_222,_GEN_223};
  assign _GEN_229 = {_GEN_226,_GEN_227};
  assign _GEN_230 = {_GEN_220,_GEN_221};
  assign _GEN_231 = {_GEN_228,_GEN_229};
  assign _GEN_232 = {_GEN_212,_GEN_213};
  assign _GEN_233 = {_GEN_230,_GEN_231};
  assign _GEN_234 = {_GEN_194,_GEN_195};
  assign _GEN_235 = {_GEN_232,_GEN_233};
  assign _GEN_236 = {_GEN_156,_GEN_157};
  assign _GEN_237 = {_GEN_234,_GEN_235};
  assign L2_meta_array_ext_RW0_wdata = {_GEN_236,_GEN_237};
endmodule
