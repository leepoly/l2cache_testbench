module TLSimpleL2Cache( // @[:freechips.rocketchip.system.DefaultConfig.fir@220955.2]
  input         clock, // @[:freechips.rocketchip.system.DefaultConfig.fir@220956.4]
  input         reset, // @[:freechips.rocketchip.system.DefaultConfig.fir@220957.4]
  output        auto_in_a_ready, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input         auto_in_a_valid, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [2:0]  auto_in_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [2:0]  auto_in_a_bits_param, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [2:0]  auto_in_a_bits_size, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [5:0]  auto_in_a_bits_source, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [32:0] auto_in_a_bits_address, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [4:0]  auto_in_a_bits_dsid, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [7:0]  auto_in_a_bits_mask, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [63:0] auto_in_a_bits_data, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input         auto_in_a_bits_corrupt, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input         auto_in_d_ready, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output        auto_in_d_valid, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [2:0]  auto_in_d_bits_opcode, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [2:0]  auto_in_d_bits_size, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [5:0]  auto_in_d_bits_source, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [63:0] auto_in_d_bits_data, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input         auto_out_a_ready, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output        auto_out_a_valid, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [2:0]  auto_out_a_bits_opcode, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [32:0] auto_out_a_bits_address, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output [63:0] auto_out_a_bits_data, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  output        auto_out_d_ready, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input         auto_out_d_valid, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [63:0] auto_out_d_bits_data, // @[:freechips.rocketchip.system.DefaultConfig.fir@220958.4]
  input  [15:0] cp_waymask, // @[:freechips.rocketchip.system.DefaultConfig.fir@220959.4]
  output [14:0] cp_capacity, // @[:freechips.rocketchip.system.DefaultConfig.fir@220959.4]
  input  [3:0]  cp_capacity_dsid // @[:freechips.rocketchip.system.DefaultConfig.fir@220959.4]
);
  wire  TLMonitor_clock; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire  TLMonitor_reset; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire  TLMonitor_io_in_a_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire  TLMonitor_io_in_a_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [2:0] TLMonitor_io_in_a_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [2:0] TLMonitor_io_in_a_bits_param; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [2:0] TLMonitor_io_in_a_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [5:0] TLMonitor_io_in_a_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [32:0] TLMonitor_io_in_a_bits_address; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [7:0] TLMonitor_io_in_a_bits_mask; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire  TLMonitor_io_in_a_bits_corrupt; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire  TLMonitor_io_in_d_ready; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire  TLMonitor_io_in_d_valid; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [2:0] TLMonitor_io_in_d_bits_opcode; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [2:0] TLMonitor_io_in_d_bits_size; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [5:0] TLMonitor_io_in_d_bits_source; // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
  wire [10:0] L2_meta_array_RW0_addr; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_en; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_clk; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wmode; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_0_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_0_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_0_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_0_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_0_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_1_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_1_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_1_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_1_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_1_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_2_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_2_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_2_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_2_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_2_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_3_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_3_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_3_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_3_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_3_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_4_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_4_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_4_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_4_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_4_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_5_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_5_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_5_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_5_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_5_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_6_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_6_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_6_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_6_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_6_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_7_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_7_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_7_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_7_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_7_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_8_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_8_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_8_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_8_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_8_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_9_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_9_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_9_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_9_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_9_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_10_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_10_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_10_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_10_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_10_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_11_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_11_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_11_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_11_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_11_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_12_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_12_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_12_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_12_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_12_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_13_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_13_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_13_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_13_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_13_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_14_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_14_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_14_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_14_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_14_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_15_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_15_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_wdata_15_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_wdata_15_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_wdata_15_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_0_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_0_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_0_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_0_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_0_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_1_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_1_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_1_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_1_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_1_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_2_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_2_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_2_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_2_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_2_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_3_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_3_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_3_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_3_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_3_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_4_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_4_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_4_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_4_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_4_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_5_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_5_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_5_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_5_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_5_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_6_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_6_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_6_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_6_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_6_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_7_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_7_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_7_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_7_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_7_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_8_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_8_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_8_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_8_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_8_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_9_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_9_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_9_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_9_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_9_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_10_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_10_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_10_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_10_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_10_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_11_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_11_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_11_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_11_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_11_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_12_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_12_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_12_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_12_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_12_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_13_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_13_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_13_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_13_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_13_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_14_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_14_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_14_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_14_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_14_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_15_valid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_15_dirty; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [15:0] L2_meta_array_RW0_rdata_15_tag; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire  L2_meta_array_RW0_rdata_15_rr_state; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [3:0] L2_meta_array_RW0_rdata_15_dsid; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
  wire [13:0] L2_data_array_RW0_addr; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_en; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_clk; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmode; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_0; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_1; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_2; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_3; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_4; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_5; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_6; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_7; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_8; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_9; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_10; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_11; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_12; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_13; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_14; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_wdata_15; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_0; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_1; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_2; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_3; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_4; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_5; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_6; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_7; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_8; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_9; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_10; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_11; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_12; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_13; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_14; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire [63:0] L2_data_array_RW0_rdata_15; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_0; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_1; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_2; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_3; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_4; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_5; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_6; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_7; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_8; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_9; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_10; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_11; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_12; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_13; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_14; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  wire  L2_data_array_RW0_wmask_15; // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
  reg [12:0] _T_258; // @[TLSimpleL2.scala 89:28:freechips.rocketchip.system.DefaultConfig.fir@221008.4]
  reg [31:0] _RAND_0;
  wire  _T_259; // @[TLSimpleL2.scala 90:26:freechips.rocketchip.system.DefaultConfig.fir@221009.4]
  wire  _T_261; // @[TLSimpleL2.scala 90:48:freechips.rocketchip.system.DefaultConfig.fir@221011.4]
  wire  _T_262; // @[TLSimpleL2.scala 90:45:freechips.rocketchip.system.DefaultConfig.fir@221012.4]
  wire [12:0] _T_264; // @[TLSimpleL2.scala 91:39:freechips.rocketchip.system.DefaultConfig.fir@221015.6]
  reg [3:0] _T_267; // @[TLSimpleL2.scala 95:22:freechips.rocketchip.system.DefaultConfig.fir@221018.4]
  reg [31:0] _RAND_1;
  wire  _T_335; // @[TLSimpleL2.scala 243:36:freechips.rocketchip.system.DefaultConfig.fir@221121.4]
  wire  _T_336; // @[TLSimpleL2.scala 243:50:freechips.rocketchip.system.DefaultConfig.fir@221122.4]
  wire  _T_337; // @[TLSimpleL2.scala 243:47:freechips.rocketchip.system.DefaultConfig.fir@221123.4]
  wire  _T_451; // @[TLSimpleL2.scala 272:45:freechips.rocketchip.system.DefaultConfig.fir@221188.4]
  wire  _T_426; // @[TLSimpleL2.scala 250:36:freechips.rocketchip.system.DefaultConfig.fir@221147.4]
  wire  _T_452; // @[TLSimpleL2.scala 272:65:freechips.rocketchip.system.DefaultConfig.fir@221189.4]
  wire  _T_273; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@221030.4]
  wire  _T_14180; // @[TLSimpleL2.scala 595:35:freechips.rocketchip.system.DefaultConfig.fir@224808.4]
  wire  _T_14199; // @[TLSimpleL2.scala 627:34:freechips.rocketchip.system.DefaultConfig.fir@224854.4]
  wire  _T_14267; // @[TLSimpleL2.scala 644:38:freechips.rocketchip.system.DefaultConfig.fir@224930.4]
  wire  _T_274; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@221033.4]
  wire  _T_275; // @[TLSimpleL2.scala 168:41:freechips.rocketchip.system.DefaultConfig.fir@221036.4]
  wire [7:0] _T_276; // @[TLSimpleL2.scala 169:45:freechips.rocketchip.system.DefaultConfig.fir@221037.4]
  wire [4:0] _T_277; // @[TLSimpleL2.scala 169:64:freechips.rocketchip.system.DefaultConfig.fir@221038.4]
  wire [5:0] _T_278; // @[TLSimpleL2.scala 169:82:freechips.rocketchip.system.DefaultConfig.fir@221039.4]
  wire [5:0] _T_279; // @[TLSimpleL2.scala 169:82:freechips.rocketchip.system.DefaultConfig.fir@221040.4]
  wire [4:0] _T_280; // @[TLSimpleL2.scala 169:82:freechips.rocketchip.system.DefaultConfig.fir@221041.4]
  wire [4:0] _T_281; // @[TLSimpleL2.scala 169:24:freechips.rocketchip.system.DefaultConfig.fir@221042.4]
  wire  _T_283; // @[TLSimpleL2.scala 174:52:freechips.rocketchip.system.DefaultConfig.fir@221044.4]
  wire  _T_284; // @[TLSimpleL2.scala 174:38:freechips.rocketchip.system.DefaultConfig.fir@221045.4]
  wire  _T_285; // @[TLSimpleL2.scala 175:53:freechips.rocketchip.system.DefaultConfig.fir@221046.4]
  wire  _T_286; // @[TLSimpleL2.scala 175:93:freechips.rocketchip.system.DefaultConfig.fir@221047.4]
  wire  _T_287; // @[TLSimpleL2.scala 175:80:freechips.rocketchip.system.DefaultConfig.fir@221048.4]
  wire  _T_288; // @[TLSimpleL2.scala 175:39:freechips.rocketchip.system.DefaultConfig.fir@221049.4]
  wire  _T_456; // @[TLSimpleL2.scala 279:31:freechips.rocketchip.system.DefaultConfig.fir@221194.4]
  wire  _T_14286; // @[TLSimpleL2.scala 664:30:freechips.rocketchip.system.DefaultConfig.fir@224952.4]
  wire  _T_14287; // @[TLSimpleL2.scala 666:33:freechips.rocketchip.system.DefaultConfig.fir@224953.4]
  wire  _T_289; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@221050.4]
  reg [32:0] _T_291; // @[TLSimpleL2.scala 182:21:freechips.rocketchip.system.DefaultConfig.fir@221051.4]
  reg [63:0] _RAND_2;
  reg [5:0] _T_293; // @[TLSimpleL2.scala 183:19:freechips.rocketchip.system.DefaultConfig.fir@221052.4]
  reg [31:0] _RAND_3;
  reg [3:0] _T_297; // @[TLSimpleL2.scala 185:25:freechips.rocketchip.system.DefaultConfig.fir@221054.4]
  reg [31:0] _RAND_4;
  reg [2:0] _T_299; // @[TLSimpleL2.scala 186:25:freechips.rocketchip.system.DefaultConfig.fir@221055.4]
  reg [31:0] _RAND_5;
  reg  _T_301; // @[TLSimpleL2.scala 188:24:freechips.rocketchip.system.DefaultConfig.fir@221056.4]
  reg [31:0] _RAND_6;
  reg  _T_303; // @[TLSimpleL2.scala 189:24:freechips.rocketchip.system.DefaultConfig.fir@221057.4]
  reg [31:0] _RAND_7;
  wire [2:0] _T_304; // @[TLSimpleL2.scala 191:31:freechips.rocketchip.system.DefaultConfig.fir@221058.4]
  reg [3:0] _T_306; // @[TLSimpleL2.scala 192:35:freechips.rocketchip.system.DefaultConfig.fir@221059.4]
  reg [31:0] _RAND_8;
  wire [4:0] _GEN_7022; // @[TLSimpleL2.scala 193:61:freechips.rocketchip.system.DefaultConfig.fir@221061.4]
  wire [4:0] _T_309; // @[TLSimpleL2.scala 193:61:freechips.rocketchip.system.DefaultConfig.fir@221062.4]
  wire [4:0] _T_310; // @[TLSimpleL2.scala 193:31:freechips.rocketchip.system.DefaultConfig.fir@221063.4]
  reg [2:0] _T_312; // @[TLSimpleL2.scala 194:41:freechips.rocketchip.system.DefaultConfig.fir@221064.4]
  reg [31:0] _RAND_9;
  wire [2:0] _T_314; // @[TLSimpleL2.scala 195:33:freechips.rocketchip.system.DefaultConfig.fir@221066.4]
  wire [4:0] _GEN_7023; // @[TLSimpleL2.scala 196:47:freechips.rocketchip.system.DefaultConfig.fir@221067.4]
  wire  _T_315; // @[TLSimpleL2.scala 196:47:freechips.rocketchip.system.DefaultConfig.fir@221067.4]
  reg [2:0] _T_317; // @[TLSimpleL2.scala 197:36:freechips.rocketchip.system.DefaultConfig.fir@221068.4]
  reg [31:0] _RAND_10;
  wire [4:0] _GEN_7024; // @[TLSimpleL2.scala 198:45:freechips.rocketchip.system.DefaultConfig.fir@221069.4]
  wire  _T_318; // @[TLSimpleL2.scala 198:45:freechips.rocketchip.system.DefaultConfig.fir@221069.4]
  reg [2:0] _T_320; // @[TLSimpleL2.scala 199:35:freechips.rocketchip.system.DefaultConfig.fir@221070.4]
  reg [31:0] _RAND_11;
  wire [4:0] _GEN_7025; // @[TLSimpleL2.scala 200:43:freechips.rocketchip.system.DefaultConfig.fir@221071.4]
  wire  _T_321; // @[TLSimpleL2.scala 200:43:freechips.rocketchip.system.DefaultConfig.fir@221071.4]
  wire [4:0] _GEN_8; // @[TLSimpleL2.scala 223:36:freechips.rocketchip.system.DefaultConfig.fir@221090.8]
  wire [4:0] _GEN_12; // @[TLSimpleL2.scala 223:36:freechips.rocketchip.system.DefaultConfig.fir@221090.8]
  wire [3:0] _GEN_13; // @[TLSimpleL2.scala 223:36:freechips.rocketchip.system.DefaultConfig.fir@221090.8]
  wire [4:0] _GEN_19; // @[TLSimpleL2.scala 207:28:freechips.rocketchip.system.DefaultConfig.fir@221074.6]
  wire [4:0] _GEN_23; // @[TLSimpleL2.scala 207:28:freechips.rocketchip.system.DefaultConfig.fir@221074.6]
  wire [3:0] _GEN_24; // @[TLSimpleL2.scala 207:28:freechips.rocketchip.system.DefaultConfig.fir@221074.6]
  wire [4:0] _GEN_30; // @[TLSimpleL2.scala 206:31:freechips.rocketchip.system.DefaultConfig.fir@221073.4]
  wire [4:0] _GEN_34; // @[TLSimpleL2.scala 206:31:freechips.rocketchip.system.DefaultConfig.fir@221073.4]
  wire [3:0] _GEN_35; // @[TLSimpleL2.scala 206:31:freechips.rocketchip.system.DefaultConfig.fir@221073.4]
  reg [63:0] _T_344_0; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_12;
  reg [63:0] _T_344_1; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_13;
  reg [63:0] _T_344_2; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_14;
  reg [63:0] _T_344_3; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_15;
  reg [63:0] _T_344_4; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_16;
  reg [63:0] _T_344_5; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_17;
  reg [63:0] _T_344_6; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_18;
  reg [63:0] _T_344_7; // @[TLSimpleL2.scala 248:29:freechips.rocketchip.system.DefaultConfig.fir@221127.4]
  reg [63:0] _RAND_19;
  reg [7:0] _T_397_0; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_20;
  reg [7:0] _T_397_1; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_21;
  reg [7:0] _T_397_2; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_22;
  reg [7:0] _T_397_3; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_23;
  reg [7:0] _T_397_4; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_24;
  reg [7:0] _T_397_5; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_25;
  reg [7:0] _T_397_6; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_26;
  reg [7:0] _T_397_7; // @[TLSimpleL2.scala 249:30:freechips.rocketchip.system.DefaultConfig.fir@221146.4]
  reg [31:0] _RAND_27;
  wire  _T_428; // @[TLSimpleL2.scala 254:60:freechips.rocketchip.system.DefaultConfig.fir@221149.4]
  wire  _T_429; // @[TLSimpleL2.scala 254:26:freechips.rocketchip.system.DefaultConfig.fir@221150.4]
  wire [2:0] _T_432; // @[TLSimpleL2.scala 256:46:freechips.rocketchip.system.DefaultConfig.fir@221155.8]
  wire [2:0] _T_435; // @[TLSimpleL2.scala 258:56:freechips.rocketchip.system.DefaultConfig.fir@221162.10]
  wire [3:0] _T_440; // @[TLSimpleL2.scala 264:56:freechips.rocketchip.system.DefaultConfig.fir@221175.6]
  wire [2:0] _T_441; // @[TLSimpleL2.scala 264:56:freechips.rocketchip.system.DefaultConfig.fir@221176.6]
  wire [3:0] _GEN_54; // @[TLSimpleL2.scala 267:33:freechips.rocketchip.system.DefaultConfig.fir@221184.6]
  wire [3:0] _GEN_72; // @[TLSimpleL2.scala 254:78:freechips.rocketchip.system.DefaultConfig.fir@221151.4]
  wire  _T_458; // @[TLSimpleL2.scala 281:36:freechips.rocketchip.system.DefaultConfig.fir@221196.4]
  wire [3:0] _GEN_73; // @[TLSimpleL2.scala 281:51:freechips.rocketchip.system.DefaultConfig.fir@221197.4]
  wire [10:0] _T_481; // @[TLSimpleL2.scala 298:21:freechips.rocketchip.system.DefaultConfig.fir@221201.4]
  wire  _T_482; // @[TLSimpleL2.scala 300:41:freechips.rocketchip.system.DefaultConfig.fir@221202.4]
  wire  _T_483; // @[TLSimpleL2.scala 300:32:freechips.rocketchip.system.DefaultConfig.fir@221203.4]
  wire  _T_484; // @[TLSimpleL2.scala 301:33:freechips.rocketchip.system.DefaultConfig.fir@221204.4]
  wire  _T_485; // @[TLSimpleL2.scala 302:61:freechips.rocketchip.system.DefaultConfig.fir@221205.4]
  wire  _T_486; // @[TLSimpleL2.scala 302:58:freechips.rocketchip.system.DefaultConfig.fir@221206.4]
  wire  _T_530_1; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221219.4]
  wire  _T_530_0; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221218.4]
  wire [1:0] _T_549; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221234.4]
  wire  _T_530_3; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221221.4]
  wire  _T_530_2; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221220.4]
  wire [1:0] _T_550; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221235.4]
  wire [3:0] _T_551; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221236.4]
  wire  _T_530_5; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221223.4]
  wire  _T_530_4; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221222.4]
  wire [1:0] _T_552; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221237.4]
  wire  _T_530_7; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221225.4]
  wire  _T_530_6; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221224.4]
  wire [1:0] _T_553; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221238.4]
  wire [3:0] _T_554; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221239.4]
  wire [7:0] _T_555; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221240.4]
  wire  _T_530_9; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221227.4]
  wire  _T_530_8; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221226.4]
  wire [1:0] _T_556; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221241.4]
  wire  _T_530_11; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221229.4]
  wire  _T_530_10; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221228.4]
  wire [1:0] _T_557; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221242.4]
  wire [3:0] _T_558; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221243.4]
  wire  _T_530_13; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221231.4]
  wire  _T_530_12; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221230.4]
  wire [1:0] _T_559; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221244.4]
  wire  _T_530_15; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221233.4]
  wire  _T_530_14; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221232.4]
  wire [1:0] _T_560; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221245.4]
  wire [3:0] _T_561; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221246.4]
  wire [7:0] _T_562; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221247.4]
  wire [15:0] _T_563; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221248.4]
  wire  _T_567_1; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221252.4]
  wire  _T_567_0; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221251.4]
  wire [1:0] _T_586; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221267.4]
  wire  _T_567_3; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221254.4]
  wire  _T_567_2; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221253.4]
  wire [1:0] _T_587; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221268.4]
  wire [3:0] _T_588; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221269.4]
  wire  _T_567_5; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221256.4]
  wire  _T_567_4; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221255.4]
  wire [1:0] _T_589; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221270.4]
  wire  _T_567_7; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221258.4]
  wire  _T_567_6; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221257.4]
  wire [1:0] _T_590; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221271.4]
  wire [3:0] _T_591; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221272.4]
  wire [7:0] _T_592; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221273.4]
  wire  _T_567_9; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221260.4]
  wire  _T_567_8; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221259.4]
  wire [1:0] _T_593; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221274.4]
  wire  _T_567_11; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221262.4]
  wire  _T_567_10; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221261.4]
  wire [1:0] _T_594; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221275.4]
  wire [3:0] _T_595; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221276.4]
  wire  _T_567_13; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221264.4]
  wire  _T_567_12; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221263.4]
  wire [1:0] _T_596; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221277.4]
  wire  _T_567_15; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221266.4]
  wire  _T_567_14; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221265.4]
  wire [1:0] _T_597; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221278.4]
  wire [3:0] _T_598; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221279.4]
  wire [7:0] _T_599; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221280.4]
  wire [15:0] _T_600; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221281.4]
  wire  _T_626_1; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221303.4]
  wire  _T_626_0; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221302.4]
  wire [1:0] _T_645; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221318.4]
  wire  _T_626_3; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221305.4]
  wire  _T_626_2; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221304.4]
  wire [1:0] _T_646; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221319.4]
  wire [3:0] _T_647; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221320.4]
  wire  _T_626_5; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221307.4]
  wire  _T_626_4; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221306.4]
  wire [1:0] _T_648; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221321.4]
  wire  _T_626_7; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221309.4]
  wire  _T_626_6; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221308.4]
  wire [1:0] _T_649; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221322.4]
  wire [3:0] _T_650; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221323.4]
  wire [7:0] _T_651; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221324.4]
  wire  _T_626_9; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221311.4]
  wire  _T_626_8; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221310.4]
  wire [1:0] _T_652; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221325.4]
  wire  _T_626_11; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221313.4]
  wire  _T_626_10; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221312.4]
  wire [1:0] _T_653; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221326.4]
  wire [3:0] _T_654; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221327.4]
  wire  _T_626_13; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221315.4]
  wire  _T_626_12; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221314.4]
  wire [1:0] _T_655; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221328.4]
  wire  _T_626_15; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221317.4]
  wire  _T_626_14; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221316.4]
  wire [1:0] _T_656; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221329.4]
  wire [3:0] _T_657; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221330.4]
  wire [7:0] _T_658; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221331.4]
  wire [15:0] _T_659; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221332.4]
  wire [3:0] _GEN_78; // @[TLSimpleL2.scala 312:39:freechips.rocketchip.system.DefaultConfig.fir@221352.4]
  reg [15:0] _T_684; // @[TLSimpleL2.scala 317:29:freechips.rocketchip.system.DefaultConfig.fir@221355.4]
  reg [31:0] _RAND_28;
  reg [15:0] _T_686; // @[TLSimpleL2.scala 318:29:freechips.rocketchip.system.DefaultConfig.fir@221356.4]
  reg [31:0] _RAND_29;
  reg [15:0] _T_690_0; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_30;
  reg [15:0] _T_690_1; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_31;
  reg [15:0] _T_690_2; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_32;
  reg [15:0] _T_690_3; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_33;
  reg [15:0] _T_690_4; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_34;
  reg [15:0] _T_690_5; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_35;
  reg [15:0] _T_690_6; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_36;
  reg [15:0] _T_690_7; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_37;
  reg [15:0] _T_690_8; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_38;
  reg [15:0] _T_690_9; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_39;
  reg [15:0] _T_690_10; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_40;
  reg [15:0] _T_690_11; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_41;
  reg [15:0] _T_690_12; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_42;
  reg [15:0] _T_690_13; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_43;
  reg [15:0] _T_690_14; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_44;
  reg [15:0] _T_690_15; // @[TLSimpleL2.scala 319:30:freechips.rocketchip.system.DefaultConfig.fir@221357.4]
  reg [31:0] _RAND_45;
  reg [15:0] _T_710; // @[TLSimpleL2.scala 320:31:freechips.rocketchip.system.DefaultConfig.fir@221358.4]
  reg [31:0] _RAND_46;
  reg [3:0] _T_714_0; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_47;
  reg [3:0] _T_714_1; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_48;
  reg [3:0] _T_714_2; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_49;
  reg [3:0] _T_714_3; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_50;
  reg [3:0] _T_714_4; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_51;
  reg [3:0] _T_714_5; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_52;
  reg [3:0] _T_714_6; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_53;
  reg [3:0] _T_714_7; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_54;
  reg [3:0] _T_714_8; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_55;
  reg [3:0] _T_714_9; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_56;
  reg [3:0] _T_714_10; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_57;
  reg [3:0] _T_714_11; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_58;
  reg [3:0] _T_714_12; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_59;
  reg [3:0] _T_714_13; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_60;
  reg [3:0] _T_714_14; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_61;
  reg [3:0] _T_714_15; // @[TLSimpleL2.scala 321:30:freechips.rocketchip.system.DefaultConfig.fir@221359.4]
  reg [31:0] _RAND_62;
  reg  _T_6887_0; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_63;
  reg  _T_6887_1; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_64;
  reg  _T_6887_2; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_65;
  reg  _T_6887_3; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_66;
  reg  _T_6887_4; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_67;
  reg  _T_6887_5; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_68;
  reg  _T_6887_6; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_69;
  reg  _T_6887_7; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_70;
  reg  _T_6887_8; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_71;
  reg  _T_6887_9; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_72;
  reg  _T_6887_10; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_73;
  reg  _T_6887_11; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_74;
  reg  _T_6887_12; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_75;
  reg  _T_6887_13; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_76;
  reg  _T_6887_14; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_77;
  reg  _T_6887_15; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_78;
  reg  _T_6887_16; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_79;
  reg  _T_6887_17; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_80;
  reg  _T_6887_18; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_81;
  reg  _T_6887_19; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_82;
  reg  _T_6887_20; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_83;
  reg  _T_6887_21; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_84;
  reg  _T_6887_22; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_85;
  reg  _T_6887_23; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_86;
  reg  _T_6887_24; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_87;
  reg  _T_6887_25; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_88;
  reg  _T_6887_26; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_89;
  reg  _T_6887_27; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_90;
  reg  _T_6887_28; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_91;
  reg  _T_6887_29; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_92;
  reg  _T_6887_30; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_93;
  reg  _T_6887_31; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_94;
  reg  _T_6887_32; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_95;
  reg  _T_6887_33; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_96;
  reg  _T_6887_34; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_97;
  reg  _T_6887_35; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_98;
  reg  _T_6887_36; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_99;
  reg  _T_6887_37; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_100;
  reg  _T_6887_38; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_101;
  reg  _T_6887_39; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_102;
  reg  _T_6887_40; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_103;
  reg  _T_6887_41; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_104;
  reg  _T_6887_42; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_105;
  reg  _T_6887_43; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_106;
  reg  _T_6887_44; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_107;
  reg  _T_6887_45; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_108;
  reg  _T_6887_46; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_109;
  reg  _T_6887_47; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_110;
  reg  _T_6887_48; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_111;
  reg  _T_6887_49; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_112;
  reg  _T_6887_50; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_113;
  reg  _T_6887_51; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_114;
  reg  _T_6887_52; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_115;
  reg  _T_6887_53; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_116;
  reg  _T_6887_54; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_117;
  reg  _T_6887_55; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_118;
  reg  _T_6887_56; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_119;
  reg  _T_6887_57; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_120;
  reg  _T_6887_58; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_121;
  reg  _T_6887_59; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_122;
  reg  _T_6887_60; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_123;
  reg  _T_6887_61; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_124;
  reg  _T_6887_62; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_125;
  reg  _T_6887_63; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_126;
  reg  _T_6887_64; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_127;
  reg  _T_6887_65; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_128;
  reg  _T_6887_66; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_129;
  reg  _T_6887_67; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_130;
  reg  _T_6887_68; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_131;
  reg  _T_6887_69; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_132;
  reg  _T_6887_70; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_133;
  reg  _T_6887_71; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_134;
  reg  _T_6887_72; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_135;
  reg  _T_6887_73; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_136;
  reg  _T_6887_74; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_137;
  reg  _T_6887_75; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_138;
  reg  _T_6887_76; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_139;
  reg  _T_6887_77; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_140;
  reg  _T_6887_78; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_141;
  reg  _T_6887_79; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_142;
  reg  _T_6887_80; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_143;
  reg  _T_6887_81; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_144;
  reg  _T_6887_82; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_145;
  reg  _T_6887_83; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_146;
  reg  _T_6887_84; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_147;
  reg  _T_6887_85; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_148;
  reg  _T_6887_86; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_149;
  reg  _T_6887_87; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_150;
  reg  _T_6887_88; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_151;
  reg  _T_6887_89; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_152;
  reg  _T_6887_90; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_153;
  reg  _T_6887_91; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_154;
  reg  _T_6887_92; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_155;
  reg  _T_6887_93; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_156;
  reg  _T_6887_94; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_157;
  reg  _T_6887_95; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_158;
  reg  _T_6887_96; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_159;
  reg  _T_6887_97; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_160;
  reg  _T_6887_98; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_161;
  reg  _T_6887_99; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_162;
  reg  _T_6887_100; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_163;
  reg  _T_6887_101; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_164;
  reg  _T_6887_102; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_165;
  reg  _T_6887_103; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_166;
  reg  _T_6887_104; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_167;
  reg  _T_6887_105; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_168;
  reg  _T_6887_106; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_169;
  reg  _T_6887_107; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_170;
  reg  _T_6887_108; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_171;
  reg  _T_6887_109; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_172;
  reg  _T_6887_110; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_173;
  reg  _T_6887_111; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_174;
  reg  _T_6887_112; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_175;
  reg  _T_6887_113; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_176;
  reg  _T_6887_114; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_177;
  reg  _T_6887_115; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_178;
  reg  _T_6887_116; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_179;
  reg  _T_6887_117; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_180;
  reg  _T_6887_118; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_181;
  reg  _T_6887_119; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_182;
  reg  _T_6887_120; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_183;
  reg  _T_6887_121; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_184;
  reg  _T_6887_122; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_185;
  reg  _T_6887_123; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_186;
  reg  _T_6887_124; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_187;
  reg  _T_6887_125; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_188;
  reg  _T_6887_126; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_189;
  reg  _T_6887_127; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_190;
  reg  _T_6887_128; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_191;
  reg  _T_6887_129; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_192;
  reg  _T_6887_130; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_193;
  reg  _T_6887_131; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_194;
  reg  _T_6887_132; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_195;
  reg  _T_6887_133; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_196;
  reg  _T_6887_134; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_197;
  reg  _T_6887_135; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_198;
  reg  _T_6887_136; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_199;
  reg  _T_6887_137; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_200;
  reg  _T_6887_138; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_201;
  reg  _T_6887_139; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_202;
  reg  _T_6887_140; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_203;
  reg  _T_6887_141; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_204;
  reg  _T_6887_142; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_205;
  reg  _T_6887_143; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_206;
  reg  _T_6887_144; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_207;
  reg  _T_6887_145; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_208;
  reg  _T_6887_146; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_209;
  reg  _T_6887_147; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_210;
  reg  _T_6887_148; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_211;
  reg  _T_6887_149; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_212;
  reg  _T_6887_150; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_213;
  reg  _T_6887_151; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_214;
  reg  _T_6887_152; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_215;
  reg  _T_6887_153; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_216;
  reg  _T_6887_154; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_217;
  reg  _T_6887_155; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_218;
  reg  _T_6887_156; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_219;
  reg  _T_6887_157; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_220;
  reg  _T_6887_158; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_221;
  reg  _T_6887_159; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_222;
  reg  _T_6887_160; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_223;
  reg  _T_6887_161; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_224;
  reg  _T_6887_162; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_225;
  reg  _T_6887_163; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_226;
  reg  _T_6887_164; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_227;
  reg  _T_6887_165; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_228;
  reg  _T_6887_166; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_229;
  reg  _T_6887_167; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_230;
  reg  _T_6887_168; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_231;
  reg  _T_6887_169; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_232;
  reg  _T_6887_170; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_233;
  reg  _T_6887_171; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_234;
  reg  _T_6887_172; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_235;
  reg  _T_6887_173; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_236;
  reg  _T_6887_174; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_237;
  reg  _T_6887_175; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_238;
  reg  _T_6887_176; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_239;
  reg  _T_6887_177; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_240;
  reg  _T_6887_178; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_241;
  reg  _T_6887_179; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_242;
  reg  _T_6887_180; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_243;
  reg  _T_6887_181; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_244;
  reg  _T_6887_182; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_245;
  reg  _T_6887_183; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_246;
  reg  _T_6887_184; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_247;
  reg  _T_6887_185; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_248;
  reg  _T_6887_186; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_249;
  reg  _T_6887_187; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_250;
  reg  _T_6887_188; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_251;
  reg  _T_6887_189; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_252;
  reg  _T_6887_190; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_253;
  reg  _T_6887_191; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_254;
  reg  _T_6887_192; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_255;
  reg  _T_6887_193; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_256;
  reg  _T_6887_194; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_257;
  reg  _T_6887_195; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_258;
  reg  _T_6887_196; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_259;
  reg  _T_6887_197; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_260;
  reg  _T_6887_198; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_261;
  reg  _T_6887_199; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_262;
  reg  _T_6887_200; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_263;
  reg  _T_6887_201; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_264;
  reg  _T_6887_202; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_265;
  reg  _T_6887_203; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_266;
  reg  _T_6887_204; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_267;
  reg  _T_6887_205; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_268;
  reg  _T_6887_206; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_269;
  reg  _T_6887_207; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_270;
  reg  _T_6887_208; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_271;
  reg  _T_6887_209; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_272;
  reg  _T_6887_210; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_273;
  reg  _T_6887_211; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_274;
  reg  _T_6887_212; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_275;
  reg  _T_6887_213; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_276;
  reg  _T_6887_214; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_277;
  reg  _T_6887_215; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_278;
  reg  _T_6887_216; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_279;
  reg  _T_6887_217; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_280;
  reg  _T_6887_218; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_281;
  reg  _T_6887_219; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_282;
  reg  _T_6887_220; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_283;
  reg  _T_6887_221; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_284;
  reg  _T_6887_222; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_285;
  reg  _T_6887_223; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_286;
  reg  _T_6887_224; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_287;
  reg  _T_6887_225; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_288;
  reg  _T_6887_226; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_289;
  reg  _T_6887_227; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_290;
  reg  _T_6887_228; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_291;
  reg  _T_6887_229; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_292;
  reg  _T_6887_230; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_293;
  reg  _T_6887_231; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_294;
  reg  _T_6887_232; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_295;
  reg  _T_6887_233; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_296;
  reg  _T_6887_234; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_297;
  reg  _T_6887_235; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_298;
  reg  _T_6887_236; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_299;
  reg  _T_6887_237; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_300;
  reg  _T_6887_238; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_301;
  reg  _T_6887_239; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_302;
  reg  _T_6887_240; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_303;
  reg  _T_6887_241; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_304;
  reg  _T_6887_242; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_305;
  reg  _T_6887_243; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_306;
  reg  _T_6887_244; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_307;
  reg  _T_6887_245; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_308;
  reg  _T_6887_246; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_309;
  reg  _T_6887_247; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_310;
  reg  _T_6887_248; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_311;
  reg  _T_6887_249; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_312;
  reg  _T_6887_250; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_313;
  reg  _T_6887_251; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_314;
  reg  _T_6887_252; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_315;
  reg  _T_6887_253; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_316;
  reg  _T_6887_254; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_317;
  reg  _T_6887_255; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_318;
  reg  _T_6887_256; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_319;
  reg  _T_6887_257; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_320;
  reg  _T_6887_258; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_321;
  reg  _T_6887_259; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_322;
  reg  _T_6887_260; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_323;
  reg  _T_6887_261; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_324;
  reg  _T_6887_262; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_325;
  reg  _T_6887_263; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_326;
  reg  _T_6887_264; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_327;
  reg  _T_6887_265; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_328;
  reg  _T_6887_266; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_329;
  reg  _T_6887_267; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_330;
  reg  _T_6887_268; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_331;
  reg  _T_6887_269; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_332;
  reg  _T_6887_270; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_333;
  reg  _T_6887_271; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_334;
  reg  _T_6887_272; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_335;
  reg  _T_6887_273; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_336;
  reg  _T_6887_274; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_337;
  reg  _T_6887_275; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_338;
  reg  _T_6887_276; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_339;
  reg  _T_6887_277; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_340;
  reg  _T_6887_278; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_341;
  reg  _T_6887_279; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_342;
  reg  _T_6887_280; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_343;
  reg  _T_6887_281; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_344;
  reg  _T_6887_282; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_345;
  reg  _T_6887_283; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_346;
  reg  _T_6887_284; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_347;
  reg  _T_6887_285; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_348;
  reg  _T_6887_286; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_349;
  reg  _T_6887_287; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_350;
  reg  _T_6887_288; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_351;
  reg  _T_6887_289; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_352;
  reg  _T_6887_290; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_353;
  reg  _T_6887_291; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_354;
  reg  _T_6887_292; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_355;
  reg  _T_6887_293; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_356;
  reg  _T_6887_294; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_357;
  reg  _T_6887_295; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_358;
  reg  _T_6887_296; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_359;
  reg  _T_6887_297; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_360;
  reg  _T_6887_298; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_361;
  reg  _T_6887_299; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_362;
  reg  _T_6887_300; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_363;
  reg  _T_6887_301; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_364;
  reg  _T_6887_302; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_365;
  reg  _T_6887_303; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_366;
  reg  _T_6887_304; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_367;
  reg  _T_6887_305; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_368;
  reg  _T_6887_306; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_369;
  reg  _T_6887_307; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_370;
  reg  _T_6887_308; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_371;
  reg  _T_6887_309; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_372;
  reg  _T_6887_310; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_373;
  reg  _T_6887_311; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_374;
  reg  _T_6887_312; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_375;
  reg  _T_6887_313; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_376;
  reg  _T_6887_314; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_377;
  reg  _T_6887_315; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_378;
  reg  _T_6887_316; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_379;
  reg  _T_6887_317; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_380;
  reg  _T_6887_318; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_381;
  reg  _T_6887_319; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_382;
  reg  _T_6887_320; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_383;
  reg  _T_6887_321; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_384;
  reg  _T_6887_322; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_385;
  reg  _T_6887_323; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_386;
  reg  _T_6887_324; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_387;
  reg  _T_6887_325; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_388;
  reg  _T_6887_326; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_389;
  reg  _T_6887_327; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_390;
  reg  _T_6887_328; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_391;
  reg  _T_6887_329; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_392;
  reg  _T_6887_330; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_393;
  reg  _T_6887_331; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_394;
  reg  _T_6887_332; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_395;
  reg  _T_6887_333; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_396;
  reg  _T_6887_334; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_397;
  reg  _T_6887_335; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_398;
  reg  _T_6887_336; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_399;
  reg  _T_6887_337; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_400;
  reg  _T_6887_338; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_401;
  reg  _T_6887_339; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_402;
  reg  _T_6887_340; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_403;
  reg  _T_6887_341; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_404;
  reg  _T_6887_342; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_405;
  reg  _T_6887_343; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_406;
  reg  _T_6887_344; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_407;
  reg  _T_6887_345; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_408;
  reg  _T_6887_346; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_409;
  reg  _T_6887_347; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_410;
  reg  _T_6887_348; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_411;
  reg  _T_6887_349; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_412;
  reg  _T_6887_350; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_413;
  reg  _T_6887_351; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_414;
  reg  _T_6887_352; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_415;
  reg  _T_6887_353; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_416;
  reg  _T_6887_354; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_417;
  reg  _T_6887_355; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_418;
  reg  _T_6887_356; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_419;
  reg  _T_6887_357; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_420;
  reg  _T_6887_358; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_421;
  reg  _T_6887_359; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_422;
  reg  _T_6887_360; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_423;
  reg  _T_6887_361; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_424;
  reg  _T_6887_362; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_425;
  reg  _T_6887_363; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_426;
  reg  _T_6887_364; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_427;
  reg  _T_6887_365; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_428;
  reg  _T_6887_366; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_429;
  reg  _T_6887_367; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_430;
  reg  _T_6887_368; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_431;
  reg  _T_6887_369; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_432;
  reg  _T_6887_370; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_433;
  reg  _T_6887_371; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_434;
  reg  _T_6887_372; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_435;
  reg  _T_6887_373; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_436;
  reg  _T_6887_374; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_437;
  reg  _T_6887_375; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_438;
  reg  _T_6887_376; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_439;
  reg  _T_6887_377; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_440;
  reg  _T_6887_378; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_441;
  reg  _T_6887_379; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_442;
  reg  _T_6887_380; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_443;
  reg  _T_6887_381; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_444;
  reg  _T_6887_382; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_445;
  reg  _T_6887_383; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_446;
  reg  _T_6887_384; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_447;
  reg  _T_6887_385; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_448;
  reg  _T_6887_386; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_449;
  reg  _T_6887_387; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_450;
  reg  _T_6887_388; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_451;
  reg  _T_6887_389; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_452;
  reg  _T_6887_390; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_453;
  reg  _T_6887_391; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_454;
  reg  _T_6887_392; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_455;
  reg  _T_6887_393; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_456;
  reg  _T_6887_394; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_457;
  reg  _T_6887_395; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_458;
  reg  _T_6887_396; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_459;
  reg  _T_6887_397; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_460;
  reg  _T_6887_398; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_461;
  reg  _T_6887_399; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_462;
  reg  _T_6887_400; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_463;
  reg  _T_6887_401; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_464;
  reg  _T_6887_402; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_465;
  reg  _T_6887_403; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_466;
  reg  _T_6887_404; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_467;
  reg  _T_6887_405; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_468;
  reg  _T_6887_406; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_469;
  reg  _T_6887_407; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_470;
  reg  _T_6887_408; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_471;
  reg  _T_6887_409; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_472;
  reg  _T_6887_410; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_473;
  reg  _T_6887_411; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_474;
  reg  _T_6887_412; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_475;
  reg  _T_6887_413; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_476;
  reg  _T_6887_414; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_477;
  reg  _T_6887_415; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_478;
  reg  _T_6887_416; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_479;
  reg  _T_6887_417; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_480;
  reg  _T_6887_418; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_481;
  reg  _T_6887_419; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_482;
  reg  _T_6887_420; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_483;
  reg  _T_6887_421; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_484;
  reg  _T_6887_422; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_485;
  reg  _T_6887_423; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_486;
  reg  _T_6887_424; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_487;
  reg  _T_6887_425; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_488;
  reg  _T_6887_426; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_489;
  reg  _T_6887_427; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_490;
  reg  _T_6887_428; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_491;
  reg  _T_6887_429; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_492;
  reg  _T_6887_430; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_493;
  reg  _T_6887_431; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_494;
  reg  _T_6887_432; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_495;
  reg  _T_6887_433; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_496;
  reg  _T_6887_434; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_497;
  reg  _T_6887_435; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_498;
  reg  _T_6887_436; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_499;
  reg  _T_6887_437; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_500;
  reg  _T_6887_438; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_501;
  reg  _T_6887_439; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_502;
  reg  _T_6887_440; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_503;
  reg  _T_6887_441; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_504;
  reg  _T_6887_442; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_505;
  reg  _T_6887_443; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_506;
  reg  _T_6887_444; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_507;
  reg  _T_6887_445; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_508;
  reg  _T_6887_446; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_509;
  reg  _T_6887_447; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_510;
  reg  _T_6887_448; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_511;
  reg  _T_6887_449; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_512;
  reg  _T_6887_450; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_513;
  reg  _T_6887_451; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_514;
  reg  _T_6887_452; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_515;
  reg  _T_6887_453; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_516;
  reg  _T_6887_454; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_517;
  reg  _T_6887_455; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_518;
  reg  _T_6887_456; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_519;
  reg  _T_6887_457; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_520;
  reg  _T_6887_458; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_521;
  reg  _T_6887_459; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_522;
  reg  _T_6887_460; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_523;
  reg  _T_6887_461; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_524;
  reg  _T_6887_462; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_525;
  reg  _T_6887_463; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_526;
  reg  _T_6887_464; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_527;
  reg  _T_6887_465; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_528;
  reg  _T_6887_466; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_529;
  reg  _T_6887_467; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_530;
  reg  _T_6887_468; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_531;
  reg  _T_6887_469; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_532;
  reg  _T_6887_470; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_533;
  reg  _T_6887_471; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_534;
  reg  _T_6887_472; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_535;
  reg  _T_6887_473; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_536;
  reg  _T_6887_474; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_537;
  reg  _T_6887_475; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_538;
  reg  _T_6887_476; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_539;
  reg  _T_6887_477; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_540;
  reg  _T_6887_478; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_541;
  reg  _T_6887_479; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_542;
  reg  _T_6887_480; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_543;
  reg  _T_6887_481; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_544;
  reg  _T_6887_482; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_545;
  reg  _T_6887_483; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_546;
  reg  _T_6887_484; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_547;
  reg  _T_6887_485; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_548;
  reg  _T_6887_486; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_549;
  reg  _T_6887_487; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_550;
  reg  _T_6887_488; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_551;
  reg  _T_6887_489; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_552;
  reg  _T_6887_490; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_553;
  reg  _T_6887_491; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_554;
  reg  _T_6887_492; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_555;
  reg  _T_6887_493; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_556;
  reg  _T_6887_494; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_557;
  reg  _T_6887_495; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_558;
  reg  _T_6887_496; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_559;
  reg  _T_6887_497; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_560;
  reg  _T_6887_498; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_561;
  reg  _T_6887_499; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_562;
  reg  _T_6887_500; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_563;
  reg  _T_6887_501; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_564;
  reg  _T_6887_502; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_565;
  reg  _T_6887_503; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_566;
  reg  _T_6887_504; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_567;
  reg  _T_6887_505; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_568;
  reg  _T_6887_506; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_569;
  reg  _T_6887_507; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_570;
  reg  _T_6887_508; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_571;
  reg  _T_6887_509; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_572;
  reg  _T_6887_510; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_573;
  reg  _T_6887_511; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_574;
  reg  _T_6887_512; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_575;
  reg  _T_6887_513; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_576;
  reg  _T_6887_514; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_577;
  reg  _T_6887_515; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_578;
  reg  _T_6887_516; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_579;
  reg  _T_6887_517; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_580;
  reg  _T_6887_518; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_581;
  reg  _T_6887_519; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_582;
  reg  _T_6887_520; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_583;
  reg  _T_6887_521; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_584;
  reg  _T_6887_522; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_585;
  reg  _T_6887_523; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_586;
  reg  _T_6887_524; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_587;
  reg  _T_6887_525; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_588;
  reg  _T_6887_526; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_589;
  reg  _T_6887_527; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_590;
  reg  _T_6887_528; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_591;
  reg  _T_6887_529; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_592;
  reg  _T_6887_530; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_593;
  reg  _T_6887_531; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_594;
  reg  _T_6887_532; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_595;
  reg  _T_6887_533; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_596;
  reg  _T_6887_534; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_597;
  reg  _T_6887_535; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_598;
  reg  _T_6887_536; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_599;
  reg  _T_6887_537; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_600;
  reg  _T_6887_538; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_601;
  reg  _T_6887_539; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_602;
  reg  _T_6887_540; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_603;
  reg  _T_6887_541; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_604;
  reg  _T_6887_542; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_605;
  reg  _T_6887_543; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_606;
  reg  _T_6887_544; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_607;
  reg  _T_6887_545; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_608;
  reg  _T_6887_546; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_609;
  reg  _T_6887_547; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_610;
  reg  _T_6887_548; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_611;
  reg  _T_6887_549; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_612;
  reg  _T_6887_550; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_613;
  reg  _T_6887_551; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_614;
  reg  _T_6887_552; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_615;
  reg  _T_6887_553; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_616;
  reg  _T_6887_554; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_617;
  reg  _T_6887_555; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_618;
  reg  _T_6887_556; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_619;
  reg  _T_6887_557; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_620;
  reg  _T_6887_558; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_621;
  reg  _T_6887_559; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_622;
  reg  _T_6887_560; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_623;
  reg  _T_6887_561; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_624;
  reg  _T_6887_562; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_625;
  reg  _T_6887_563; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_626;
  reg  _T_6887_564; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_627;
  reg  _T_6887_565; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_628;
  reg  _T_6887_566; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_629;
  reg  _T_6887_567; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_630;
  reg  _T_6887_568; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_631;
  reg  _T_6887_569; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_632;
  reg  _T_6887_570; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_633;
  reg  _T_6887_571; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_634;
  reg  _T_6887_572; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_635;
  reg  _T_6887_573; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_636;
  reg  _T_6887_574; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_637;
  reg  _T_6887_575; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_638;
  reg  _T_6887_576; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_639;
  reg  _T_6887_577; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_640;
  reg  _T_6887_578; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_641;
  reg  _T_6887_579; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_642;
  reg  _T_6887_580; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_643;
  reg  _T_6887_581; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_644;
  reg  _T_6887_582; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_645;
  reg  _T_6887_583; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_646;
  reg  _T_6887_584; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_647;
  reg  _T_6887_585; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_648;
  reg  _T_6887_586; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_649;
  reg  _T_6887_587; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_650;
  reg  _T_6887_588; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_651;
  reg  _T_6887_589; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_652;
  reg  _T_6887_590; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_653;
  reg  _T_6887_591; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_654;
  reg  _T_6887_592; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_655;
  reg  _T_6887_593; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_656;
  reg  _T_6887_594; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_657;
  reg  _T_6887_595; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_658;
  reg  _T_6887_596; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_659;
  reg  _T_6887_597; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_660;
  reg  _T_6887_598; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_661;
  reg  _T_6887_599; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_662;
  reg  _T_6887_600; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_663;
  reg  _T_6887_601; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_664;
  reg  _T_6887_602; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_665;
  reg  _T_6887_603; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_666;
  reg  _T_6887_604; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_667;
  reg  _T_6887_605; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_668;
  reg  _T_6887_606; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_669;
  reg  _T_6887_607; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_670;
  reg  _T_6887_608; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_671;
  reg  _T_6887_609; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_672;
  reg  _T_6887_610; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_673;
  reg  _T_6887_611; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_674;
  reg  _T_6887_612; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_675;
  reg  _T_6887_613; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_676;
  reg  _T_6887_614; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_677;
  reg  _T_6887_615; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_678;
  reg  _T_6887_616; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_679;
  reg  _T_6887_617; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_680;
  reg  _T_6887_618; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_681;
  reg  _T_6887_619; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_682;
  reg  _T_6887_620; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_683;
  reg  _T_6887_621; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_684;
  reg  _T_6887_622; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_685;
  reg  _T_6887_623; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_686;
  reg  _T_6887_624; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_687;
  reg  _T_6887_625; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_688;
  reg  _T_6887_626; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_689;
  reg  _T_6887_627; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_690;
  reg  _T_6887_628; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_691;
  reg  _T_6887_629; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_692;
  reg  _T_6887_630; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_693;
  reg  _T_6887_631; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_694;
  reg  _T_6887_632; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_695;
  reg  _T_6887_633; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_696;
  reg  _T_6887_634; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_697;
  reg  _T_6887_635; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_698;
  reg  _T_6887_636; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_699;
  reg  _T_6887_637; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_700;
  reg  _T_6887_638; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_701;
  reg  _T_6887_639; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_702;
  reg  _T_6887_640; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_703;
  reg  _T_6887_641; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_704;
  reg  _T_6887_642; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_705;
  reg  _T_6887_643; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_706;
  reg  _T_6887_644; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_707;
  reg  _T_6887_645; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_708;
  reg  _T_6887_646; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_709;
  reg  _T_6887_647; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_710;
  reg  _T_6887_648; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_711;
  reg  _T_6887_649; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_712;
  reg  _T_6887_650; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_713;
  reg  _T_6887_651; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_714;
  reg  _T_6887_652; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_715;
  reg  _T_6887_653; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_716;
  reg  _T_6887_654; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_717;
  reg  _T_6887_655; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_718;
  reg  _T_6887_656; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_719;
  reg  _T_6887_657; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_720;
  reg  _T_6887_658; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_721;
  reg  _T_6887_659; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_722;
  reg  _T_6887_660; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_723;
  reg  _T_6887_661; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_724;
  reg  _T_6887_662; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_725;
  reg  _T_6887_663; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_726;
  reg  _T_6887_664; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_727;
  reg  _T_6887_665; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_728;
  reg  _T_6887_666; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_729;
  reg  _T_6887_667; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_730;
  reg  _T_6887_668; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_731;
  reg  _T_6887_669; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_732;
  reg  _T_6887_670; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_733;
  reg  _T_6887_671; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_734;
  reg  _T_6887_672; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_735;
  reg  _T_6887_673; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_736;
  reg  _T_6887_674; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_737;
  reg  _T_6887_675; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_738;
  reg  _T_6887_676; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_739;
  reg  _T_6887_677; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_740;
  reg  _T_6887_678; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_741;
  reg  _T_6887_679; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_742;
  reg  _T_6887_680; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_743;
  reg  _T_6887_681; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_744;
  reg  _T_6887_682; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_745;
  reg  _T_6887_683; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_746;
  reg  _T_6887_684; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_747;
  reg  _T_6887_685; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_748;
  reg  _T_6887_686; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_749;
  reg  _T_6887_687; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_750;
  reg  _T_6887_688; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_751;
  reg  _T_6887_689; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_752;
  reg  _T_6887_690; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_753;
  reg  _T_6887_691; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_754;
  reg  _T_6887_692; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_755;
  reg  _T_6887_693; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_756;
  reg  _T_6887_694; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_757;
  reg  _T_6887_695; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_758;
  reg  _T_6887_696; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_759;
  reg  _T_6887_697; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_760;
  reg  _T_6887_698; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_761;
  reg  _T_6887_699; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_762;
  reg  _T_6887_700; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_763;
  reg  _T_6887_701; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_764;
  reg  _T_6887_702; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_765;
  reg  _T_6887_703; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_766;
  reg  _T_6887_704; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_767;
  reg  _T_6887_705; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_768;
  reg  _T_6887_706; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_769;
  reg  _T_6887_707; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_770;
  reg  _T_6887_708; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_771;
  reg  _T_6887_709; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_772;
  reg  _T_6887_710; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_773;
  reg  _T_6887_711; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_774;
  reg  _T_6887_712; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_775;
  reg  _T_6887_713; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_776;
  reg  _T_6887_714; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_777;
  reg  _T_6887_715; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_778;
  reg  _T_6887_716; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_779;
  reg  _T_6887_717; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_780;
  reg  _T_6887_718; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_781;
  reg  _T_6887_719; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_782;
  reg  _T_6887_720; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_783;
  reg  _T_6887_721; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_784;
  reg  _T_6887_722; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_785;
  reg  _T_6887_723; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_786;
  reg  _T_6887_724; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_787;
  reg  _T_6887_725; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_788;
  reg  _T_6887_726; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_789;
  reg  _T_6887_727; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_790;
  reg  _T_6887_728; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_791;
  reg  _T_6887_729; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_792;
  reg  _T_6887_730; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_793;
  reg  _T_6887_731; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_794;
  reg  _T_6887_732; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_795;
  reg  _T_6887_733; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_796;
  reg  _T_6887_734; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_797;
  reg  _T_6887_735; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_798;
  reg  _T_6887_736; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_799;
  reg  _T_6887_737; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_800;
  reg  _T_6887_738; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_801;
  reg  _T_6887_739; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_802;
  reg  _T_6887_740; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_803;
  reg  _T_6887_741; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_804;
  reg  _T_6887_742; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_805;
  reg  _T_6887_743; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_806;
  reg  _T_6887_744; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_807;
  reg  _T_6887_745; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_808;
  reg  _T_6887_746; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_809;
  reg  _T_6887_747; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_810;
  reg  _T_6887_748; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_811;
  reg  _T_6887_749; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_812;
  reg  _T_6887_750; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_813;
  reg  _T_6887_751; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_814;
  reg  _T_6887_752; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_815;
  reg  _T_6887_753; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_816;
  reg  _T_6887_754; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_817;
  reg  _T_6887_755; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_818;
  reg  _T_6887_756; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_819;
  reg  _T_6887_757; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_820;
  reg  _T_6887_758; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_821;
  reg  _T_6887_759; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_822;
  reg  _T_6887_760; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_823;
  reg  _T_6887_761; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_824;
  reg  _T_6887_762; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_825;
  reg  _T_6887_763; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_826;
  reg  _T_6887_764; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_827;
  reg  _T_6887_765; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_828;
  reg  _T_6887_766; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_829;
  reg  _T_6887_767; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_830;
  reg  _T_6887_768; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_831;
  reg  _T_6887_769; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_832;
  reg  _T_6887_770; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_833;
  reg  _T_6887_771; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_834;
  reg  _T_6887_772; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_835;
  reg  _T_6887_773; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_836;
  reg  _T_6887_774; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_837;
  reg  _T_6887_775; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_838;
  reg  _T_6887_776; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_839;
  reg  _T_6887_777; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_840;
  reg  _T_6887_778; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_841;
  reg  _T_6887_779; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_842;
  reg  _T_6887_780; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_843;
  reg  _T_6887_781; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_844;
  reg  _T_6887_782; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_845;
  reg  _T_6887_783; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_846;
  reg  _T_6887_784; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_847;
  reg  _T_6887_785; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_848;
  reg  _T_6887_786; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_849;
  reg  _T_6887_787; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_850;
  reg  _T_6887_788; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_851;
  reg  _T_6887_789; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_852;
  reg  _T_6887_790; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_853;
  reg  _T_6887_791; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_854;
  reg  _T_6887_792; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_855;
  reg  _T_6887_793; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_856;
  reg  _T_6887_794; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_857;
  reg  _T_6887_795; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_858;
  reg  _T_6887_796; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_859;
  reg  _T_6887_797; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_860;
  reg  _T_6887_798; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_861;
  reg  _T_6887_799; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_862;
  reg  _T_6887_800; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_863;
  reg  _T_6887_801; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_864;
  reg  _T_6887_802; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_865;
  reg  _T_6887_803; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_866;
  reg  _T_6887_804; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_867;
  reg  _T_6887_805; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_868;
  reg  _T_6887_806; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_869;
  reg  _T_6887_807; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_870;
  reg  _T_6887_808; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_871;
  reg  _T_6887_809; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_872;
  reg  _T_6887_810; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_873;
  reg  _T_6887_811; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_874;
  reg  _T_6887_812; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_875;
  reg  _T_6887_813; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_876;
  reg  _T_6887_814; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_877;
  reg  _T_6887_815; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_878;
  reg  _T_6887_816; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_879;
  reg  _T_6887_817; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_880;
  reg  _T_6887_818; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_881;
  reg  _T_6887_819; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_882;
  reg  _T_6887_820; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_883;
  reg  _T_6887_821; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_884;
  reg  _T_6887_822; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_885;
  reg  _T_6887_823; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_886;
  reg  _T_6887_824; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_887;
  reg  _T_6887_825; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_888;
  reg  _T_6887_826; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_889;
  reg  _T_6887_827; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_890;
  reg  _T_6887_828; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_891;
  reg  _T_6887_829; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_892;
  reg  _T_6887_830; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_893;
  reg  _T_6887_831; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_894;
  reg  _T_6887_832; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_895;
  reg  _T_6887_833; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_896;
  reg  _T_6887_834; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_897;
  reg  _T_6887_835; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_898;
  reg  _T_6887_836; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_899;
  reg  _T_6887_837; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_900;
  reg  _T_6887_838; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_901;
  reg  _T_6887_839; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_902;
  reg  _T_6887_840; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_903;
  reg  _T_6887_841; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_904;
  reg  _T_6887_842; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_905;
  reg  _T_6887_843; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_906;
  reg  _T_6887_844; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_907;
  reg  _T_6887_845; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_908;
  reg  _T_6887_846; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_909;
  reg  _T_6887_847; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_910;
  reg  _T_6887_848; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_911;
  reg  _T_6887_849; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_912;
  reg  _T_6887_850; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_913;
  reg  _T_6887_851; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_914;
  reg  _T_6887_852; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_915;
  reg  _T_6887_853; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_916;
  reg  _T_6887_854; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_917;
  reg  _T_6887_855; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_918;
  reg  _T_6887_856; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_919;
  reg  _T_6887_857; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_920;
  reg  _T_6887_858; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_921;
  reg  _T_6887_859; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_922;
  reg  _T_6887_860; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_923;
  reg  _T_6887_861; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_924;
  reg  _T_6887_862; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_925;
  reg  _T_6887_863; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_926;
  reg  _T_6887_864; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_927;
  reg  _T_6887_865; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_928;
  reg  _T_6887_866; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_929;
  reg  _T_6887_867; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_930;
  reg  _T_6887_868; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_931;
  reg  _T_6887_869; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_932;
  reg  _T_6887_870; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_933;
  reg  _T_6887_871; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_934;
  reg  _T_6887_872; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_935;
  reg  _T_6887_873; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_936;
  reg  _T_6887_874; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_937;
  reg  _T_6887_875; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_938;
  reg  _T_6887_876; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_939;
  reg  _T_6887_877; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_940;
  reg  _T_6887_878; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_941;
  reg  _T_6887_879; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_942;
  reg  _T_6887_880; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_943;
  reg  _T_6887_881; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_944;
  reg  _T_6887_882; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_945;
  reg  _T_6887_883; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_946;
  reg  _T_6887_884; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_947;
  reg  _T_6887_885; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_948;
  reg  _T_6887_886; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_949;
  reg  _T_6887_887; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_950;
  reg  _T_6887_888; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_951;
  reg  _T_6887_889; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_952;
  reg  _T_6887_890; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_953;
  reg  _T_6887_891; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_954;
  reg  _T_6887_892; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_955;
  reg  _T_6887_893; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_956;
  reg  _T_6887_894; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_957;
  reg  _T_6887_895; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_958;
  reg  _T_6887_896; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_959;
  reg  _T_6887_897; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_960;
  reg  _T_6887_898; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_961;
  reg  _T_6887_899; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_962;
  reg  _T_6887_900; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_963;
  reg  _T_6887_901; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_964;
  reg  _T_6887_902; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_965;
  reg  _T_6887_903; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_966;
  reg  _T_6887_904; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_967;
  reg  _T_6887_905; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_968;
  reg  _T_6887_906; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_969;
  reg  _T_6887_907; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_970;
  reg  _T_6887_908; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_971;
  reg  _T_6887_909; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_972;
  reg  _T_6887_910; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_973;
  reg  _T_6887_911; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_974;
  reg  _T_6887_912; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_975;
  reg  _T_6887_913; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_976;
  reg  _T_6887_914; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_977;
  reg  _T_6887_915; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_978;
  reg  _T_6887_916; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_979;
  reg  _T_6887_917; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_980;
  reg  _T_6887_918; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_981;
  reg  _T_6887_919; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_982;
  reg  _T_6887_920; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_983;
  reg  _T_6887_921; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_984;
  reg  _T_6887_922; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_985;
  reg  _T_6887_923; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_986;
  reg  _T_6887_924; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_987;
  reg  _T_6887_925; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_988;
  reg  _T_6887_926; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_989;
  reg  _T_6887_927; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_990;
  reg  _T_6887_928; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_991;
  reg  _T_6887_929; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_992;
  reg  _T_6887_930; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_993;
  reg  _T_6887_931; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_994;
  reg  _T_6887_932; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_995;
  reg  _T_6887_933; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_996;
  reg  _T_6887_934; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_997;
  reg  _T_6887_935; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_998;
  reg  _T_6887_936; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_999;
  reg  _T_6887_937; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1000;
  reg  _T_6887_938; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1001;
  reg  _T_6887_939; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1002;
  reg  _T_6887_940; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1003;
  reg  _T_6887_941; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1004;
  reg  _T_6887_942; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1005;
  reg  _T_6887_943; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1006;
  reg  _T_6887_944; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1007;
  reg  _T_6887_945; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1008;
  reg  _T_6887_946; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1009;
  reg  _T_6887_947; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1010;
  reg  _T_6887_948; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1011;
  reg  _T_6887_949; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1012;
  reg  _T_6887_950; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1013;
  reg  _T_6887_951; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1014;
  reg  _T_6887_952; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1015;
  reg  _T_6887_953; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1016;
  reg  _T_6887_954; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1017;
  reg  _T_6887_955; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1018;
  reg  _T_6887_956; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1019;
  reg  _T_6887_957; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1020;
  reg  _T_6887_958; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1021;
  reg  _T_6887_959; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1022;
  reg  _T_6887_960; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1023;
  reg  _T_6887_961; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1024;
  reg  _T_6887_962; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1025;
  reg  _T_6887_963; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1026;
  reg  _T_6887_964; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1027;
  reg  _T_6887_965; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1028;
  reg  _T_6887_966; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1029;
  reg  _T_6887_967; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1030;
  reg  _T_6887_968; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1031;
  reg  _T_6887_969; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1032;
  reg  _T_6887_970; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1033;
  reg  _T_6887_971; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1034;
  reg  _T_6887_972; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1035;
  reg  _T_6887_973; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1036;
  reg  _T_6887_974; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1037;
  reg  _T_6887_975; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1038;
  reg  _T_6887_976; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1039;
  reg  _T_6887_977; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1040;
  reg  _T_6887_978; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1041;
  reg  _T_6887_979; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1042;
  reg  _T_6887_980; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1043;
  reg  _T_6887_981; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1044;
  reg  _T_6887_982; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1045;
  reg  _T_6887_983; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1046;
  reg  _T_6887_984; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1047;
  reg  _T_6887_985; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1048;
  reg  _T_6887_986; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1049;
  reg  _T_6887_987; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1050;
  reg  _T_6887_988; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1051;
  reg  _T_6887_989; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1052;
  reg  _T_6887_990; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1053;
  reg  _T_6887_991; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1054;
  reg  _T_6887_992; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1055;
  reg  _T_6887_993; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1056;
  reg  _T_6887_994; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1057;
  reg  _T_6887_995; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1058;
  reg  _T_6887_996; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1059;
  reg  _T_6887_997; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1060;
  reg  _T_6887_998; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1061;
  reg  _T_6887_999; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1062;
  reg  _T_6887_1000; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1063;
  reg  _T_6887_1001; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1064;
  reg  _T_6887_1002; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1065;
  reg  _T_6887_1003; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1066;
  reg  _T_6887_1004; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1067;
  reg  _T_6887_1005; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1068;
  reg  _T_6887_1006; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1069;
  reg  _T_6887_1007; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1070;
  reg  _T_6887_1008; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1071;
  reg  _T_6887_1009; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1072;
  reg  _T_6887_1010; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1073;
  reg  _T_6887_1011; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1074;
  reg  _T_6887_1012; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1075;
  reg  _T_6887_1013; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1076;
  reg  _T_6887_1014; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1077;
  reg  _T_6887_1015; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1078;
  reg  _T_6887_1016; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1079;
  reg  _T_6887_1017; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1080;
  reg  _T_6887_1018; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1081;
  reg  _T_6887_1019; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1082;
  reg  _T_6887_1020; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1083;
  reg  _T_6887_1021; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1084;
  reg  _T_6887_1022; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1085;
  reg  _T_6887_1023; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1086;
  reg  _T_6887_1024; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1087;
  reg  _T_6887_1025; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1088;
  reg  _T_6887_1026; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1089;
  reg  _T_6887_1027; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1090;
  reg  _T_6887_1028; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1091;
  reg  _T_6887_1029; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1092;
  reg  _T_6887_1030; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1093;
  reg  _T_6887_1031; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1094;
  reg  _T_6887_1032; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1095;
  reg  _T_6887_1033; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1096;
  reg  _T_6887_1034; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1097;
  reg  _T_6887_1035; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1098;
  reg  _T_6887_1036; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1099;
  reg  _T_6887_1037; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1100;
  reg  _T_6887_1038; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1101;
  reg  _T_6887_1039; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1102;
  reg  _T_6887_1040; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1103;
  reg  _T_6887_1041; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1104;
  reg  _T_6887_1042; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1105;
  reg  _T_6887_1043; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1106;
  reg  _T_6887_1044; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1107;
  reg  _T_6887_1045; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1108;
  reg  _T_6887_1046; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1109;
  reg  _T_6887_1047; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1110;
  reg  _T_6887_1048; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1111;
  reg  _T_6887_1049; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1112;
  reg  _T_6887_1050; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1113;
  reg  _T_6887_1051; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1114;
  reg  _T_6887_1052; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1115;
  reg  _T_6887_1053; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1116;
  reg  _T_6887_1054; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1117;
  reg  _T_6887_1055; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1118;
  reg  _T_6887_1056; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1119;
  reg  _T_6887_1057; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1120;
  reg  _T_6887_1058; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1121;
  reg  _T_6887_1059; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1122;
  reg  _T_6887_1060; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1123;
  reg  _T_6887_1061; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1124;
  reg  _T_6887_1062; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1125;
  reg  _T_6887_1063; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1126;
  reg  _T_6887_1064; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1127;
  reg  _T_6887_1065; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1128;
  reg  _T_6887_1066; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1129;
  reg  _T_6887_1067; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1130;
  reg  _T_6887_1068; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1131;
  reg  _T_6887_1069; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1132;
  reg  _T_6887_1070; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1133;
  reg  _T_6887_1071; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1134;
  reg  _T_6887_1072; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1135;
  reg  _T_6887_1073; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1136;
  reg  _T_6887_1074; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1137;
  reg  _T_6887_1075; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1138;
  reg  _T_6887_1076; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1139;
  reg  _T_6887_1077; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1140;
  reg  _T_6887_1078; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1141;
  reg  _T_6887_1079; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1142;
  reg  _T_6887_1080; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1143;
  reg  _T_6887_1081; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1144;
  reg  _T_6887_1082; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1145;
  reg  _T_6887_1083; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1146;
  reg  _T_6887_1084; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1147;
  reg  _T_6887_1085; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1148;
  reg  _T_6887_1086; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1149;
  reg  _T_6887_1087; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1150;
  reg  _T_6887_1088; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1151;
  reg  _T_6887_1089; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1152;
  reg  _T_6887_1090; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1153;
  reg  _T_6887_1091; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1154;
  reg  _T_6887_1092; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1155;
  reg  _T_6887_1093; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1156;
  reg  _T_6887_1094; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1157;
  reg  _T_6887_1095; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1158;
  reg  _T_6887_1096; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1159;
  reg  _T_6887_1097; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1160;
  reg  _T_6887_1098; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1161;
  reg  _T_6887_1099; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1162;
  reg  _T_6887_1100; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1163;
  reg  _T_6887_1101; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1164;
  reg  _T_6887_1102; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1165;
  reg  _T_6887_1103; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1166;
  reg  _T_6887_1104; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1167;
  reg  _T_6887_1105; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1168;
  reg  _T_6887_1106; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1169;
  reg  _T_6887_1107; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1170;
  reg  _T_6887_1108; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1171;
  reg  _T_6887_1109; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1172;
  reg  _T_6887_1110; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1173;
  reg  _T_6887_1111; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1174;
  reg  _T_6887_1112; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1175;
  reg  _T_6887_1113; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1176;
  reg  _T_6887_1114; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1177;
  reg  _T_6887_1115; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1178;
  reg  _T_6887_1116; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1179;
  reg  _T_6887_1117; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1180;
  reg  _T_6887_1118; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1181;
  reg  _T_6887_1119; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1182;
  reg  _T_6887_1120; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1183;
  reg  _T_6887_1121; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1184;
  reg  _T_6887_1122; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1185;
  reg  _T_6887_1123; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1186;
  reg  _T_6887_1124; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1187;
  reg  _T_6887_1125; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1188;
  reg  _T_6887_1126; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1189;
  reg  _T_6887_1127; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1190;
  reg  _T_6887_1128; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1191;
  reg  _T_6887_1129; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1192;
  reg  _T_6887_1130; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1193;
  reg  _T_6887_1131; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1194;
  reg  _T_6887_1132; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1195;
  reg  _T_6887_1133; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1196;
  reg  _T_6887_1134; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1197;
  reg  _T_6887_1135; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1198;
  reg  _T_6887_1136; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1199;
  reg  _T_6887_1137; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1200;
  reg  _T_6887_1138; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1201;
  reg  _T_6887_1139; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1202;
  reg  _T_6887_1140; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1203;
  reg  _T_6887_1141; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1204;
  reg  _T_6887_1142; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1205;
  reg  _T_6887_1143; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1206;
  reg  _T_6887_1144; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1207;
  reg  _T_6887_1145; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1208;
  reg  _T_6887_1146; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1209;
  reg  _T_6887_1147; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1210;
  reg  _T_6887_1148; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1211;
  reg  _T_6887_1149; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1212;
  reg  _T_6887_1150; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1213;
  reg  _T_6887_1151; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1214;
  reg  _T_6887_1152; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1215;
  reg  _T_6887_1153; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1216;
  reg  _T_6887_1154; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1217;
  reg  _T_6887_1155; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1218;
  reg  _T_6887_1156; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1219;
  reg  _T_6887_1157; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1220;
  reg  _T_6887_1158; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1221;
  reg  _T_6887_1159; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1222;
  reg  _T_6887_1160; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1223;
  reg  _T_6887_1161; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1224;
  reg  _T_6887_1162; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1225;
  reg  _T_6887_1163; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1226;
  reg  _T_6887_1164; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1227;
  reg  _T_6887_1165; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1228;
  reg  _T_6887_1166; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1229;
  reg  _T_6887_1167; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1230;
  reg  _T_6887_1168; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1231;
  reg  _T_6887_1169; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1232;
  reg  _T_6887_1170; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1233;
  reg  _T_6887_1171; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1234;
  reg  _T_6887_1172; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1235;
  reg  _T_6887_1173; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1236;
  reg  _T_6887_1174; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1237;
  reg  _T_6887_1175; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1238;
  reg  _T_6887_1176; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1239;
  reg  _T_6887_1177; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1240;
  reg  _T_6887_1178; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1241;
  reg  _T_6887_1179; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1242;
  reg  _T_6887_1180; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1243;
  reg  _T_6887_1181; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1244;
  reg  _T_6887_1182; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1245;
  reg  _T_6887_1183; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1246;
  reg  _T_6887_1184; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1247;
  reg  _T_6887_1185; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1248;
  reg  _T_6887_1186; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1249;
  reg  _T_6887_1187; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1250;
  reg  _T_6887_1188; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1251;
  reg  _T_6887_1189; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1252;
  reg  _T_6887_1190; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1253;
  reg  _T_6887_1191; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1254;
  reg  _T_6887_1192; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1255;
  reg  _T_6887_1193; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1256;
  reg  _T_6887_1194; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1257;
  reg  _T_6887_1195; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1258;
  reg  _T_6887_1196; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1259;
  reg  _T_6887_1197; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1260;
  reg  _T_6887_1198; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1261;
  reg  _T_6887_1199; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1262;
  reg  _T_6887_1200; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1263;
  reg  _T_6887_1201; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1264;
  reg  _T_6887_1202; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1265;
  reg  _T_6887_1203; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1266;
  reg  _T_6887_1204; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1267;
  reg  _T_6887_1205; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1268;
  reg  _T_6887_1206; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1269;
  reg  _T_6887_1207; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1270;
  reg  _T_6887_1208; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1271;
  reg  _T_6887_1209; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1272;
  reg  _T_6887_1210; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1273;
  reg  _T_6887_1211; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1274;
  reg  _T_6887_1212; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1275;
  reg  _T_6887_1213; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1276;
  reg  _T_6887_1214; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1277;
  reg  _T_6887_1215; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1278;
  reg  _T_6887_1216; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1279;
  reg  _T_6887_1217; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1280;
  reg  _T_6887_1218; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1281;
  reg  _T_6887_1219; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1282;
  reg  _T_6887_1220; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1283;
  reg  _T_6887_1221; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1284;
  reg  _T_6887_1222; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1285;
  reg  _T_6887_1223; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1286;
  reg  _T_6887_1224; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1287;
  reg  _T_6887_1225; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1288;
  reg  _T_6887_1226; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1289;
  reg  _T_6887_1227; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1290;
  reg  _T_6887_1228; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1291;
  reg  _T_6887_1229; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1292;
  reg  _T_6887_1230; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1293;
  reg  _T_6887_1231; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1294;
  reg  _T_6887_1232; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1295;
  reg  _T_6887_1233; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1296;
  reg  _T_6887_1234; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1297;
  reg  _T_6887_1235; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1298;
  reg  _T_6887_1236; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1299;
  reg  _T_6887_1237; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1300;
  reg  _T_6887_1238; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1301;
  reg  _T_6887_1239; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1302;
  reg  _T_6887_1240; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1303;
  reg  _T_6887_1241; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1304;
  reg  _T_6887_1242; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1305;
  reg  _T_6887_1243; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1306;
  reg  _T_6887_1244; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1307;
  reg  _T_6887_1245; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1308;
  reg  _T_6887_1246; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1309;
  reg  _T_6887_1247; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1310;
  reg  _T_6887_1248; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1311;
  reg  _T_6887_1249; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1312;
  reg  _T_6887_1250; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1313;
  reg  _T_6887_1251; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1314;
  reg  _T_6887_1252; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1315;
  reg  _T_6887_1253; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1316;
  reg  _T_6887_1254; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1317;
  reg  _T_6887_1255; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1318;
  reg  _T_6887_1256; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1319;
  reg  _T_6887_1257; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1320;
  reg  _T_6887_1258; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1321;
  reg  _T_6887_1259; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1322;
  reg  _T_6887_1260; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1323;
  reg  _T_6887_1261; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1324;
  reg  _T_6887_1262; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1325;
  reg  _T_6887_1263; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1326;
  reg  _T_6887_1264; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1327;
  reg  _T_6887_1265; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1328;
  reg  _T_6887_1266; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1329;
  reg  _T_6887_1267; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1330;
  reg  _T_6887_1268; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1331;
  reg  _T_6887_1269; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1332;
  reg  _T_6887_1270; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1333;
  reg  _T_6887_1271; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1334;
  reg  _T_6887_1272; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1335;
  reg  _T_6887_1273; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1336;
  reg  _T_6887_1274; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1337;
  reg  _T_6887_1275; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1338;
  reg  _T_6887_1276; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1339;
  reg  _T_6887_1277; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1340;
  reg  _T_6887_1278; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1341;
  reg  _T_6887_1279; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1342;
  reg  _T_6887_1280; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1343;
  reg  _T_6887_1281; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1344;
  reg  _T_6887_1282; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1345;
  reg  _T_6887_1283; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1346;
  reg  _T_6887_1284; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1347;
  reg  _T_6887_1285; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1348;
  reg  _T_6887_1286; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1349;
  reg  _T_6887_1287; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1350;
  reg  _T_6887_1288; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1351;
  reg  _T_6887_1289; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1352;
  reg  _T_6887_1290; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1353;
  reg  _T_6887_1291; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1354;
  reg  _T_6887_1292; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1355;
  reg  _T_6887_1293; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1356;
  reg  _T_6887_1294; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1357;
  reg  _T_6887_1295; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1358;
  reg  _T_6887_1296; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1359;
  reg  _T_6887_1297; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1360;
  reg  _T_6887_1298; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1361;
  reg  _T_6887_1299; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1362;
  reg  _T_6887_1300; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1363;
  reg  _T_6887_1301; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1364;
  reg  _T_6887_1302; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1365;
  reg  _T_6887_1303; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1366;
  reg  _T_6887_1304; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1367;
  reg  _T_6887_1305; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1368;
  reg  _T_6887_1306; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1369;
  reg  _T_6887_1307; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1370;
  reg  _T_6887_1308; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1371;
  reg  _T_6887_1309; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1372;
  reg  _T_6887_1310; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1373;
  reg  _T_6887_1311; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1374;
  reg  _T_6887_1312; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1375;
  reg  _T_6887_1313; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1376;
  reg  _T_6887_1314; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1377;
  reg  _T_6887_1315; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1378;
  reg  _T_6887_1316; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1379;
  reg  _T_6887_1317; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1380;
  reg  _T_6887_1318; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1381;
  reg  _T_6887_1319; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1382;
  reg  _T_6887_1320; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1383;
  reg  _T_6887_1321; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1384;
  reg  _T_6887_1322; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1385;
  reg  _T_6887_1323; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1386;
  reg  _T_6887_1324; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1387;
  reg  _T_6887_1325; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1388;
  reg  _T_6887_1326; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1389;
  reg  _T_6887_1327; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1390;
  reg  _T_6887_1328; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1391;
  reg  _T_6887_1329; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1392;
  reg  _T_6887_1330; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1393;
  reg  _T_6887_1331; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1394;
  reg  _T_6887_1332; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1395;
  reg  _T_6887_1333; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1396;
  reg  _T_6887_1334; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1397;
  reg  _T_6887_1335; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1398;
  reg  _T_6887_1336; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1399;
  reg  _T_6887_1337; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1400;
  reg  _T_6887_1338; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1401;
  reg  _T_6887_1339; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1402;
  reg  _T_6887_1340; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1403;
  reg  _T_6887_1341; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1404;
  reg  _T_6887_1342; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1405;
  reg  _T_6887_1343; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1406;
  reg  _T_6887_1344; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1407;
  reg  _T_6887_1345; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1408;
  reg  _T_6887_1346; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1409;
  reg  _T_6887_1347; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1410;
  reg  _T_6887_1348; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1411;
  reg  _T_6887_1349; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1412;
  reg  _T_6887_1350; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1413;
  reg  _T_6887_1351; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1414;
  reg  _T_6887_1352; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1415;
  reg  _T_6887_1353; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1416;
  reg  _T_6887_1354; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1417;
  reg  _T_6887_1355; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1418;
  reg  _T_6887_1356; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1419;
  reg  _T_6887_1357; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1420;
  reg  _T_6887_1358; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1421;
  reg  _T_6887_1359; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1422;
  reg  _T_6887_1360; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1423;
  reg  _T_6887_1361; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1424;
  reg  _T_6887_1362; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1425;
  reg  _T_6887_1363; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1426;
  reg  _T_6887_1364; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1427;
  reg  _T_6887_1365; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1428;
  reg  _T_6887_1366; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1429;
  reg  _T_6887_1367; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1430;
  reg  _T_6887_1368; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1431;
  reg  _T_6887_1369; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1432;
  reg  _T_6887_1370; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1433;
  reg  _T_6887_1371; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1434;
  reg  _T_6887_1372; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1435;
  reg  _T_6887_1373; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1436;
  reg  _T_6887_1374; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1437;
  reg  _T_6887_1375; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1438;
  reg  _T_6887_1376; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1439;
  reg  _T_6887_1377; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1440;
  reg  _T_6887_1378; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1441;
  reg  _T_6887_1379; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1442;
  reg  _T_6887_1380; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1443;
  reg  _T_6887_1381; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1444;
  reg  _T_6887_1382; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1445;
  reg  _T_6887_1383; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1446;
  reg  _T_6887_1384; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1447;
  reg  _T_6887_1385; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1448;
  reg  _T_6887_1386; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1449;
  reg  _T_6887_1387; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1450;
  reg  _T_6887_1388; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1451;
  reg  _T_6887_1389; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1452;
  reg  _T_6887_1390; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1453;
  reg  _T_6887_1391; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1454;
  reg  _T_6887_1392; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1455;
  reg  _T_6887_1393; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1456;
  reg  _T_6887_1394; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1457;
  reg  _T_6887_1395; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1458;
  reg  _T_6887_1396; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1459;
  reg  _T_6887_1397; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1460;
  reg  _T_6887_1398; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1461;
  reg  _T_6887_1399; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1462;
  reg  _T_6887_1400; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1463;
  reg  _T_6887_1401; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1464;
  reg  _T_6887_1402; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1465;
  reg  _T_6887_1403; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1466;
  reg  _T_6887_1404; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1467;
  reg  _T_6887_1405; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1468;
  reg  _T_6887_1406; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1469;
  reg  _T_6887_1407; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1470;
  reg  _T_6887_1408; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1471;
  reg  _T_6887_1409; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1472;
  reg  _T_6887_1410; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1473;
  reg  _T_6887_1411; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1474;
  reg  _T_6887_1412; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1475;
  reg  _T_6887_1413; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1476;
  reg  _T_6887_1414; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1477;
  reg  _T_6887_1415; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1478;
  reg  _T_6887_1416; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1479;
  reg  _T_6887_1417; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1480;
  reg  _T_6887_1418; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1481;
  reg  _T_6887_1419; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1482;
  reg  _T_6887_1420; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1483;
  reg  _T_6887_1421; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1484;
  reg  _T_6887_1422; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1485;
  reg  _T_6887_1423; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1486;
  reg  _T_6887_1424; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1487;
  reg  _T_6887_1425; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1488;
  reg  _T_6887_1426; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1489;
  reg  _T_6887_1427; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1490;
  reg  _T_6887_1428; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1491;
  reg  _T_6887_1429; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1492;
  reg  _T_6887_1430; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1493;
  reg  _T_6887_1431; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1494;
  reg  _T_6887_1432; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1495;
  reg  _T_6887_1433; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1496;
  reg  _T_6887_1434; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1497;
  reg  _T_6887_1435; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1498;
  reg  _T_6887_1436; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1499;
  reg  _T_6887_1437; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1500;
  reg  _T_6887_1438; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1501;
  reg  _T_6887_1439; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1502;
  reg  _T_6887_1440; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1503;
  reg  _T_6887_1441; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1504;
  reg  _T_6887_1442; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1505;
  reg  _T_6887_1443; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1506;
  reg  _T_6887_1444; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1507;
  reg  _T_6887_1445; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1508;
  reg  _T_6887_1446; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1509;
  reg  _T_6887_1447; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1510;
  reg  _T_6887_1448; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1511;
  reg  _T_6887_1449; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1512;
  reg  _T_6887_1450; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1513;
  reg  _T_6887_1451; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1514;
  reg  _T_6887_1452; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1515;
  reg  _T_6887_1453; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1516;
  reg  _T_6887_1454; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1517;
  reg  _T_6887_1455; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1518;
  reg  _T_6887_1456; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1519;
  reg  _T_6887_1457; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1520;
  reg  _T_6887_1458; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1521;
  reg  _T_6887_1459; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1522;
  reg  _T_6887_1460; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1523;
  reg  _T_6887_1461; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1524;
  reg  _T_6887_1462; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1525;
  reg  _T_6887_1463; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1526;
  reg  _T_6887_1464; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1527;
  reg  _T_6887_1465; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1528;
  reg  _T_6887_1466; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1529;
  reg  _T_6887_1467; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1530;
  reg  _T_6887_1468; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1531;
  reg  _T_6887_1469; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1532;
  reg  _T_6887_1470; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1533;
  reg  _T_6887_1471; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1534;
  reg  _T_6887_1472; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1535;
  reg  _T_6887_1473; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1536;
  reg  _T_6887_1474; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1537;
  reg  _T_6887_1475; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1538;
  reg  _T_6887_1476; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1539;
  reg  _T_6887_1477; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1540;
  reg  _T_6887_1478; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1541;
  reg  _T_6887_1479; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1542;
  reg  _T_6887_1480; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1543;
  reg  _T_6887_1481; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1544;
  reg  _T_6887_1482; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1545;
  reg  _T_6887_1483; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1546;
  reg  _T_6887_1484; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1547;
  reg  _T_6887_1485; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1548;
  reg  _T_6887_1486; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1549;
  reg  _T_6887_1487; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1550;
  reg  _T_6887_1488; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1551;
  reg  _T_6887_1489; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1552;
  reg  _T_6887_1490; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1553;
  reg  _T_6887_1491; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1554;
  reg  _T_6887_1492; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1555;
  reg  _T_6887_1493; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1556;
  reg  _T_6887_1494; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1557;
  reg  _T_6887_1495; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1558;
  reg  _T_6887_1496; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1559;
  reg  _T_6887_1497; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1560;
  reg  _T_6887_1498; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1561;
  reg  _T_6887_1499; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1562;
  reg  _T_6887_1500; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1563;
  reg  _T_6887_1501; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1564;
  reg  _T_6887_1502; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1565;
  reg  _T_6887_1503; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1566;
  reg  _T_6887_1504; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1567;
  reg  _T_6887_1505; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1568;
  reg  _T_6887_1506; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1569;
  reg  _T_6887_1507; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1570;
  reg  _T_6887_1508; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1571;
  reg  _T_6887_1509; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1572;
  reg  _T_6887_1510; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1573;
  reg  _T_6887_1511; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1574;
  reg  _T_6887_1512; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1575;
  reg  _T_6887_1513; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1576;
  reg  _T_6887_1514; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1577;
  reg  _T_6887_1515; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1578;
  reg  _T_6887_1516; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1579;
  reg  _T_6887_1517; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1580;
  reg  _T_6887_1518; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1581;
  reg  _T_6887_1519; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1582;
  reg  _T_6887_1520; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1583;
  reg  _T_6887_1521; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1584;
  reg  _T_6887_1522; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1585;
  reg  _T_6887_1523; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1586;
  reg  _T_6887_1524; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1587;
  reg  _T_6887_1525; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1588;
  reg  _T_6887_1526; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1589;
  reg  _T_6887_1527; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1590;
  reg  _T_6887_1528; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1591;
  reg  _T_6887_1529; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1592;
  reg  _T_6887_1530; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1593;
  reg  _T_6887_1531; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1594;
  reg  _T_6887_1532; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1595;
  reg  _T_6887_1533; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1596;
  reg  _T_6887_1534; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1597;
  reg  _T_6887_1535; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1598;
  reg  _T_6887_1536; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1599;
  reg  _T_6887_1537; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1600;
  reg  _T_6887_1538; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1601;
  reg  _T_6887_1539; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1602;
  reg  _T_6887_1540; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1603;
  reg  _T_6887_1541; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1604;
  reg  _T_6887_1542; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1605;
  reg  _T_6887_1543; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1606;
  reg  _T_6887_1544; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1607;
  reg  _T_6887_1545; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1608;
  reg  _T_6887_1546; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1609;
  reg  _T_6887_1547; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1610;
  reg  _T_6887_1548; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1611;
  reg  _T_6887_1549; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1612;
  reg  _T_6887_1550; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1613;
  reg  _T_6887_1551; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1614;
  reg  _T_6887_1552; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1615;
  reg  _T_6887_1553; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1616;
  reg  _T_6887_1554; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1617;
  reg  _T_6887_1555; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1618;
  reg  _T_6887_1556; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1619;
  reg  _T_6887_1557; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1620;
  reg  _T_6887_1558; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1621;
  reg  _T_6887_1559; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1622;
  reg  _T_6887_1560; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1623;
  reg  _T_6887_1561; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1624;
  reg  _T_6887_1562; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1625;
  reg  _T_6887_1563; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1626;
  reg  _T_6887_1564; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1627;
  reg  _T_6887_1565; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1628;
  reg  _T_6887_1566; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1629;
  reg  _T_6887_1567; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1630;
  reg  _T_6887_1568; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1631;
  reg  _T_6887_1569; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1632;
  reg  _T_6887_1570; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1633;
  reg  _T_6887_1571; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1634;
  reg  _T_6887_1572; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1635;
  reg  _T_6887_1573; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1636;
  reg  _T_6887_1574; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1637;
  reg  _T_6887_1575; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1638;
  reg  _T_6887_1576; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1639;
  reg  _T_6887_1577; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1640;
  reg  _T_6887_1578; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1641;
  reg  _T_6887_1579; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1642;
  reg  _T_6887_1580; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1643;
  reg  _T_6887_1581; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1644;
  reg  _T_6887_1582; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1645;
  reg  _T_6887_1583; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1646;
  reg  _T_6887_1584; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1647;
  reg  _T_6887_1585; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1648;
  reg  _T_6887_1586; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1649;
  reg  _T_6887_1587; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1650;
  reg  _T_6887_1588; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1651;
  reg  _T_6887_1589; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1652;
  reg  _T_6887_1590; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1653;
  reg  _T_6887_1591; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1654;
  reg  _T_6887_1592; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1655;
  reg  _T_6887_1593; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1656;
  reg  _T_6887_1594; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1657;
  reg  _T_6887_1595; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1658;
  reg  _T_6887_1596; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1659;
  reg  _T_6887_1597; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1660;
  reg  _T_6887_1598; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1661;
  reg  _T_6887_1599; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1662;
  reg  _T_6887_1600; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1663;
  reg  _T_6887_1601; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1664;
  reg  _T_6887_1602; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1665;
  reg  _T_6887_1603; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1666;
  reg  _T_6887_1604; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1667;
  reg  _T_6887_1605; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1668;
  reg  _T_6887_1606; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1669;
  reg  _T_6887_1607; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1670;
  reg  _T_6887_1608; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1671;
  reg  _T_6887_1609; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1672;
  reg  _T_6887_1610; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1673;
  reg  _T_6887_1611; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1674;
  reg  _T_6887_1612; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1675;
  reg  _T_6887_1613; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1676;
  reg  _T_6887_1614; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1677;
  reg  _T_6887_1615; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1678;
  reg  _T_6887_1616; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1679;
  reg  _T_6887_1617; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1680;
  reg  _T_6887_1618; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1681;
  reg  _T_6887_1619; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1682;
  reg  _T_6887_1620; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1683;
  reg  _T_6887_1621; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1684;
  reg  _T_6887_1622; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1685;
  reg  _T_6887_1623; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1686;
  reg  _T_6887_1624; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1687;
  reg  _T_6887_1625; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1688;
  reg  _T_6887_1626; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1689;
  reg  _T_6887_1627; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1690;
  reg  _T_6887_1628; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1691;
  reg  _T_6887_1629; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1692;
  reg  _T_6887_1630; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1693;
  reg  _T_6887_1631; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1694;
  reg  _T_6887_1632; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1695;
  reg  _T_6887_1633; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1696;
  reg  _T_6887_1634; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1697;
  reg  _T_6887_1635; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1698;
  reg  _T_6887_1636; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1699;
  reg  _T_6887_1637; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1700;
  reg  _T_6887_1638; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1701;
  reg  _T_6887_1639; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1702;
  reg  _T_6887_1640; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1703;
  reg  _T_6887_1641; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1704;
  reg  _T_6887_1642; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1705;
  reg  _T_6887_1643; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1706;
  reg  _T_6887_1644; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1707;
  reg  _T_6887_1645; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1708;
  reg  _T_6887_1646; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1709;
  reg  _T_6887_1647; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1710;
  reg  _T_6887_1648; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1711;
  reg  _T_6887_1649; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1712;
  reg  _T_6887_1650; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1713;
  reg  _T_6887_1651; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1714;
  reg  _T_6887_1652; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1715;
  reg  _T_6887_1653; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1716;
  reg  _T_6887_1654; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1717;
  reg  _T_6887_1655; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1718;
  reg  _T_6887_1656; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1719;
  reg  _T_6887_1657; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1720;
  reg  _T_6887_1658; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1721;
  reg  _T_6887_1659; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1722;
  reg  _T_6887_1660; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1723;
  reg  _T_6887_1661; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1724;
  reg  _T_6887_1662; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1725;
  reg  _T_6887_1663; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1726;
  reg  _T_6887_1664; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1727;
  reg  _T_6887_1665; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1728;
  reg  _T_6887_1666; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1729;
  reg  _T_6887_1667; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1730;
  reg  _T_6887_1668; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1731;
  reg  _T_6887_1669; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1732;
  reg  _T_6887_1670; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1733;
  reg  _T_6887_1671; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1734;
  reg  _T_6887_1672; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1735;
  reg  _T_6887_1673; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1736;
  reg  _T_6887_1674; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1737;
  reg  _T_6887_1675; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1738;
  reg  _T_6887_1676; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1739;
  reg  _T_6887_1677; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1740;
  reg  _T_6887_1678; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1741;
  reg  _T_6887_1679; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1742;
  reg  _T_6887_1680; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1743;
  reg  _T_6887_1681; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1744;
  reg  _T_6887_1682; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1745;
  reg  _T_6887_1683; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1746;
  reg  _T_6887_1684; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1747;
  reg  _T_6887_1685; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1748;
  reg  _T_6887_1686; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1749;
  reg  _T_6887_1687; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1750;
  reg  _T_6887_1688; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1751;
  reg  _T_6887_1689; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1752;
  reg  _T_6887_1690; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1753;
  reg  _T_6887_1691; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1754;
  reg  _T_6887_1692; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1755;
  reg  _T_6887_1693; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1756;
  reg  _T_6887_1694; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1757;
  reg  _T_6887_1695; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1758;
  reg  _T_6887_1696; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1759;
  reg  _T_6887_1697; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1760;
  reg  _T_6887_1698; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1761;
  reg  _T_6887_1699; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1762;
  reg  _T_6887_1700; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1763;
  reg  _T_6887_1701; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1764;
  reg  _T_6887_1702; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1765;
  reg  _T_6887_1703; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1766;
  reg  _T_6887_1704; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1767;
  reg  _T_6887_1705; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1768;
  reg  _T_6887_1706; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1769;
  reg  _T_6887_1707; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1770;
  reg  _T_6887_1708; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1771;
  reg  _T_6887_1709; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1772;
  reg  _T_6887_1710; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1773;
  reg  _T_6887_1711; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1774;
  reg  _T_6887_1712; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1775;
  reg  _T_6887_1713; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1776;
  reg  _T_6887_1714; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1777;
  reg  _T_6887_1715; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1778;
  reg  _T_6887_1716; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1779;
  reg  _T_6887_1717; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1780;
  reg  _T_6887_1718; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1781;
  reg  _T_6887_1719; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1782;
  reg  _T_6887_1720; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1783;
  reg  _T_6887_1721; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1784;
  reg  _T_6887_1722; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1785;
  reg  _T_6887_1723; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1786;
  reg  _T_6887_1724; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1787;
  reg  _T_6887_1725; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1788;
  reg  _T_6887_1726; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1789;
  reg  _T_6887_1727; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1790;
  reg  _T_6887_1728; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1791;
  reg  _T_6887_1729; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1792;
  reg  _T_6887_1730; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1793;
  reg  _T_6887_1731; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1794;
  reg  _T_6887_1732; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1795;
  reg  _T_6887_1733; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1796;
  reg  _T_6887_1734; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1797;
  reg  _T_6887_1735; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1798;
  reg  _T_6887_1736; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1799;
  reg  _T_6887_1737; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1800;
  reg  _T_6887_1738; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1801;
  reg  _T_6887_1739; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1802;
  reg  _T_6887_1740; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1803;
  reg  _T_6887_1741; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1804;
  reg  _T_6887_1742; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1805;
  reg  _T_6887_1743; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1806;
  reg  _T_6887_1744; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1807;
  reg  _T_6887_1745; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1808;
  reg  _T_6887_1746; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1809;
  reg  _T_6887_1747; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1810;
  reg  _T_6887_1748; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1811;
  reg  _T_6887_1749; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1812;
  reg  _T_6887_1750; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1813;
  reg  _T_6887_1751; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1814;
  reg  _T_6887_1752; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1815;
  reg  _T_6887_1753; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1816;
  reg  _T_6887_1754; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1817;
  reg  _T_6887_1755; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1818;
  reg  _T_6887_1756; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1819;
  reg  _T_6887_1757; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1820;
  reg  _T_6887_1758; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1821;
  reg  _T_6887_1759; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1822;
  reg  _T_6887_1760; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1823;
  reg  _T_6887_1761; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1824;
  reg  _T_6887_1762; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1825;
  reg  _T_6887_1763; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1826;
  reg  _T_6887_1764; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1827;
  reg  _T_6887_1765; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1828;
  reg  _T_6887_1766; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1829;
  reg  _T_6887_1767; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1830;
  reg  _T_6887_1768; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1831;
  reg  _T_6887_1769; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1832;
  reg  _T_6887_1770; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1833;
  reg  _T_6887_1771; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1834;
  reg  _T_6887_1772; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1835;
  reg  _T_6887_1773; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1836;
  reg  _T_6887_1774; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1837;
  reg  _T_6887_1775; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1838;
  reg  _T_6887_1776; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1839;
  reg  _T_6887_1777; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1840;
  reg  _T_6887_1778; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1841;
  reg  _T_6887_1779; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1842;
  reg  _T_6887_1780; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1843;
  reg  _T_6887_1781; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1844;
  reg  _T_6887_1782; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1845;
  reg  _T_6887_1783; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1846;
  reg  _T_6887_1784; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1847;
  reg  _T_6887_1785; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1848;
  reg  _T_6887_1786; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1849;
  reg  _T_6887_1787; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1850;
  reg  _T_6887_1788; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1851;
  reg  _T_6887_1789; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1852;
  reg  _T_6887_1790; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1853;
  reg  _T_6887_1791; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1854;
  reg  _T_6887_1792; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1855;
  reg  _T_6887_1793; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1856;
  reg  _T_6887_1794; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1857;
  reg  _T_6887_1795; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1858;
  reg  _T_6887_1796; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1859;
  reg  _T_6887_1797; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1860;
  reg  _T_6887_1798; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1861;
  reg  _T_6887_1799; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1862;
  reg  _T_6887_1800; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1863;
  reg  _T_6887_1801; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1864;
  reg  _T_6887_1802; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1865;
  reg  _T_6887_1803; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1866;
  reg  _T_6887_1804; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1867;
  reg  _T_6887_1805; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1868;
  reg  _T_6887_1806; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1869;
  reg  _T_6887_1807; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1870;
  reg  _T_6887_1808; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1871;
  reg  _T_6887_1809; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1872;
  reg  _T_6887_1810; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1873;
  reg  _T_6887_1811; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1874;
  reg  _T_6887_1812; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1875;
  reg  _T_6887_1813; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1876;
  reg  _T_6887_1814; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1877;
  reg  _T_6887_1815; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1878;
  reg  _T_6887_1816; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1879;
  reg  _T_6887_1817; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1880;
  reg  _T_6887_1818; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1881;
  reg  _T_6887_1819; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1882;
  reg  _T_6887_1820; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1883;
  reg  _T_6887_1821; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1884;
  reg  _T_6887_1822; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1885;
  reg  _T_6887_1823; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1886;
  reg  _T_6887_1824; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1887;
  reg  _T_6887_1825; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1888;
  reg  _T_6887_1826; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1889;
  reg  _T_6887_1827; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1890;
  reg  _T_6887_1828; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1891;
  reg  _T_6887_1829; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1892;
  reg  _T_6887_1830; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1893;
  reg  _T_6887_1831; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1894;
  reg  _T_6887_1832; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1895;
  reg  _T_6887_1833; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1896;
  reg  _T_6887_1834; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1897;
  reg  _T_6887_1835; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1898;
  reg  _T_6887_1836; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1899;
  reg  _T_6887_1837; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1900;
  reg  _T_6887_1838; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1901;
  reg  _T_6887_1839; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1902;
  reg  _T_6887_1840; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1903;
  reg  _T_6887_1841; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1904;
  reg  _T_6887_1842; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1905;
  reg  _T_6887_1843; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1906;
  reg  _T_6887_1844; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1907;
  reg  _T_6887_1845; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1908;
  reg  _T_6887_1846; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1909;
  reg  _T_6887_1847; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1910;
  reg  _T_6887_1848; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1911;
  reg  _T_6887_1849; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1912;
  reg  _T_6887_1850; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1913;
  reg  _T_6887_1851; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1914;
  reg  _T_6887_1852; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1915;
  reg  _T_6887_1853; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1916;
  reg  _T_6887_1854; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1917;
  reg  _T_6887_1855; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1918;
  reg  _T_6887_1856; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1919;
  reg  _T_6887_1857; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1920;
  reg  _T_6887_1858; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1921;
  reg  _T_6887_1859; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1922;
  reg  _T_6887_1860; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1923;
  reg  _T_6887_1861; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1924;
  reg  _T_6887_1862; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1925;
  reg  _T_6887_1863; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1926;
  reg  _T_6887_1864; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1927;
  reg  _T_6887_1865; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1928;
  reg  _T_6887_1866; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1929;
  reg  _T_6887_1867; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1930;
  reg  _T_6887_1868; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1931;
  reg  _T_6887_1869; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1932;
  reg  _T_6887_1870; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1933;
  reg  _T_6887_1871; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1934;
  reg  _T_6887_1872; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1935;
  reg  _T_6887_1873; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1936;
  reg  _T_6887_1874; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1937;
  reg  _T_6887_1875; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1938;
  reg  _T_6887_1876; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1939;
  reg  _T_6887_1877; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1940;
  reg  _T_6887_1878; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1941;
  reg  _T_6887_1879; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1942;
  reg  _T_6887_1880; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1943;
  reg  _T_6887_1881; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1944;
  reg  _T_6887_1882; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1945;
  reg  _T_6887_1883; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1946;
  reg  _T_6887_1884; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1947;
  reg  _T_6887_1885; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1948;
  reg  _T_6887_1886; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1949;
  reg  _T_6887_1887; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1950;
  reg  _T_6887_1888; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1951;
  reg  _T_6887_1889; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1952;
  reg  _T_6887_1890; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1953;
  reg  _T_6887_1891; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1954;
  reg  _T_6887_1892; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1955;
  reg  _T_6887_1893; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1956;
  reg  _T_6887_1894; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1957;
  reg  _T_6887_1895; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1958;
  reg  _T_6887_1896; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1959;
  reg  _T_6887_1897; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1960;
  reg  _T_6887_1898; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1961;
  reg  _T_6887_1899; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1962;
  reg  _T_6887_1900; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1963;
  reg  _T_6887_1901; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1964;
  reg  _T_6887_1902; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1965;
  reg  _T_6887_1903; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1966;
  reg  _T_6887_1904; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1967;
  reg  _T_6887_1905; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1968;
  reg  _T_6887_1906; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1969;
  reg  _T_6887_1907; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1970;
  reg  _T_6887_1908; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1971;
  reg  _T_6887_1909; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1972;
  reg  _T_6887_1910; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1973;
  reg  _T_6887_1911; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1974;
  reg  _T_6887_1912; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1975;
  reg  _T_6887_1913; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1976;
  reg  _T_6887_1914; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1977;
  reg  _T_6887_1915; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1978;
  reg  _T_6887_1916; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1979;
  reg  _T_6887_1917; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1980;
  reg  _T_6887_1918; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1981;
  reg  _T_6887_1919; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1982;
  reg  _T_6887_1920; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1983;
  reg  _T_6887_1921; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1984;
  reg  _T_6887_1922; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1985;
  reg  _T_6887_1923; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1986;
  reg  _T_6887_1924; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1987;
  reg  _T_6887_1925; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1988;
  reg  _T_6887_1926; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1989;
  reg  _T_6887_1927; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1990;
  reg  _T_6887_1928; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1991;
  reg  _T_6887_1929; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1992;
  reg  _T_6887_1930; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1993;
  reg  _T_6887_1931; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1994;
  reg  _T_6887_1932; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1995;
  reg  _T_6887_1933; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1996;
  reg  _T_6887_1934; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1997;
  reg  _T_6887_1935; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1998;
  reg  _T_6887_1936; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_1999;
  reg  _T_6887_1937; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2000;
  reg  _T_6887_1938; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2001;
  reg  _T_6887_1939; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2002;
  reg  _T_6887_1940; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2003;
  reg  _T_6887_1941; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2004;
  reg  _T_6887_1942; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2005;
  reg  _T_6887_1943; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2006;
  reg  _T_6887_1944; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2007;
  reg  _T_6887_1945; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2008;
  reg  _T_6887_1946; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2009;
  reg  _T_6887_1947; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2010;
  reg  _T_6887_1948; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2011;
  reg  _T_6887_1949; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2012;
  reg  _T_6887_1950; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2013;
  reg  _T_6887_1951; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2014;
  reg  _T_6887_1952; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2015;
  reg  _T_6887_1953; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2016;
  reg  _T_6887_1954; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2017;
  reg  _T_6887_1955; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2018;
  reg  _T_6887_1956; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2019;
  reg  _T_6887_1957; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2020;
  reg  _T_6887_1958; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2021;
  reg  _T_6887_1959; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2022;
  reg  _T_6887_1960; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2023;
  reg  _T_6887_1961; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2024;
  reg  _T_6887_1962; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2025;
  reg  _T_6887_1963; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2026;
  reg  _T_6887_1964; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2027;
  reg  _T_6887_1965; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2028;
  reg  _T_6887_1966; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2029;
  reg  _T_6887_1967; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2030;
  reg  _T_6887_1968; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2031;
  reg  _T_6887_1969; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2032;
  reg  _T_6887_1970; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2033;
  reg  _T_6887_1971; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2034;
  reg  _T_6887_1972; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2035;
  reg  _T_6887_1973; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2036;
  reg  _T_6887_1974; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2037;
  reg  _T_6887_1975; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2038;
  reg  _T_6887_1976; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2039;
  reg  _T_6887_1977; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2040;
  reg  _T_6887_1978; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2041;
  reg  _T_6887_1979; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2042;
  reg  _T_6887_1980; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2043;
  reg  _T_6887_1981; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2044;
  reg  _T_6887_1982; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2045;
  reg  _T_6887_1983; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2046;
  reg  _T_6887_1984; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2047;
  reg  _T_6887_1985; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2048;
  reg  _T_6887_1986; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2049;
  reg  _T_6887_1987; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2050;
  reg  _T_6887_1988; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2051;
  reg  _T_6887_1989; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2052;
  reg  _T_6887_1990; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2053;
  reg  _T_6887_1991; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2054;
  reg  _T_6887_1992; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2055;
  reg  _T_6887_1993; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2056;
  reg  _T_6887_1994; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2057;
  reg  _T_6887_1995; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2058;
  reg  _T_6887_1996; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2059;
  reg  _T_6887_1997; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2060;
  reg  _T_6887_1998; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2061;
  reg  _T_6887_1999; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2062;
  reg  _T_6887_2000; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2063;
  reg  _T_6887_2001; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2064;
  reg  _T_6887_2002; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2065;
  reg  _T_6887_2003; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2066;
  reg  _T_6887_2004; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2067;
  reg  _T_6887_2005; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2068;
  reg  _T_6887_2006; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2069;
  reg  _T_6887_2007; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2070;
  reg  _T_6887_2008; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2071;
  reg  _T_6887_2009; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2072;
  reg  _T_6887_2010; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2073;
  reg  _T_6887_2011; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2074;
  reg  _T_6887_2012; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2075;
  reg  _T_6887_2013; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2076;
  reg  _T_6887_2014; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2077;
  reg  _T_6887_2015; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2078;
  reg  _T_6887_2016; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2079;
  reg  _T_6887_2017; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2080;
  reg  _T_6887_2018; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2081;
  reg  _T_6887_2019; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2082;
  reg  _T_6887_2020; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2083;
  reg  _T_6887_2021; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2084;
  reg  _T_6887_2022; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2085;
  reg  _T_6887_2023; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2086;
  reg  _T_6887_2024; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2087;
  reg  _T_6887_2025; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2088;
  reg  _T_6887_2026; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2089;
  reg  _T_6887_2027; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2090;
  reg  _T_6887_2028; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2091;
  reg  _T_6887_2029; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2092;
  reg  _T_6887_2030; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2093;
  reg  _T_6887_2031; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2094;
  reg  _T_6887_2032; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2095;
  reg  _T_6887_2033; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2096;
  reg  _T_6887_2034; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2097;
  reg  _T_6887_2035; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2098;
  reg  _T_6887_2036; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2099;
  reg  _T_6887_2037; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2100;
  reg  _T_6887_2038; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2101;
  reg  _T_6887_2039; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2102;
  reg  _T_6887_2040; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2103;
  reg  _T_6887_2041; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2104;
  reg  _T_6887_2042; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2105;
  reg  _T_6887_2043; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2106;
  reg  _T_6887_2044; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2107;
  reg  _T_6887_2045; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2108;
  reg  _T_6887_2046; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2109;
  reg  _T_6887_2047; // @[TLSimpleL2.scala 323:42:freechips.rocketchip.system.DefaultConfig.fir@223410.4]
  reg [31:0] _RAND_2110;
  wire  _T_13036; // @[TLSimpleL2.scala 326:19:freechips.rocketchip.system.DefaultConfig.fir@223411.4]
  wire  _GEN_80; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_81; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_82; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_83; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_84; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_85; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_86; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_87; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_88; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_89; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_90; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_91; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_92; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_93; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_94; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_95; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_96; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_97; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_98; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_99; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_100; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_101; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_102; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_103; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_104; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_105; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_106; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_107; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_108; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_109; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_110; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_111; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_112; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_113; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_114; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_115; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_116; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_117; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_118; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_119; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_120; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_121; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_122; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_123; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_124; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_125; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_126; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_127; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_128; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_129; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_130; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_131; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_132; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_133; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_134; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_135; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_136; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_137; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_138; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_139; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_140; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_141; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_142; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_143; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_144; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_145; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_146; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_147; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_148; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_149; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_150; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_151; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_152; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_153; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_154; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_155; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_156; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_157; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_158; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_159; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_160; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_161; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_162; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_163; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_164; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_165; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_166; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_167; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_168; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_169; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_170; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_171; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_172; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_173; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_174; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_175; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_176; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_177; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_178; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_179; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_180; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_181; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_182; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_183; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_184; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_185; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_186; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_187; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_188; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_189; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_190; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_191; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_192; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_193; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_194; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_195; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_196; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_197; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_198; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_199; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_200; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_201; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_202; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_203; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_204; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_205; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_206; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_207; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_208; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_209; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_210; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_211; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_212; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_213; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_214; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_215; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_216; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_217; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_218; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_219; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_220; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_221; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_222; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_223; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_224; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_225; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_226; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_227; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_228; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_229; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_230; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_231; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_232; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_233; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_234; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_235; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_236; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_237; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_238; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_239; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_240; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_241; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_242; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_243; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_244; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_245; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_246; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_247; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_248; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_249; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_250; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_251; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_252; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_253; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_254; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_255; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_256; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_257; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_258; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_259; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_260; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_261; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_262; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_263; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_264; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_265; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_266; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_267; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_268; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_269; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_270; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_271; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_272; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_273; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_274; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_275; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_276; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_277; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_278; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_279; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_280; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_281; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_282; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_283; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_284; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_285; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_286; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_287; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_288; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_289; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_290; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_291; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_292; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_293; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_294; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_295; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_296; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_297; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_298; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_299; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_300; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_301; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_302; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_303; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_304; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_305; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_306; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_307; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_308; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_309; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_310; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_311; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_312; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_313; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_314; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_315; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_316; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_317; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_318; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_319; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_320; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_321; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_322; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_323; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_324; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_325; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_326; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_327; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_328; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_329; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_330; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_331; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_332; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_333; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_334; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_335; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_336; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_337; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_338; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_339; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_340; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_341; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_342; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_343; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_344; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_345; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_346; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_347; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_348; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_349; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_350; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_351; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_352; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_353; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_354; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_355; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_356; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_357; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_358; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_359; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_360; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_361; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_362; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_363; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_364; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_365; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_366; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_367; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_368; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_369; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_370; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_371; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_372; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_373; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_374; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_375; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_376; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_377; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_378; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_379; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_380; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_381; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_382; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_383; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_384; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_385; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_386; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_387; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_388; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_389; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_390; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_391; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_392; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_393; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_394; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_395; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_396; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_397; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_398; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_399; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_400; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_401; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_402; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_403; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_404; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_405; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_406; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_407; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_408; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_409; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_410; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_411; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_412; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_413; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_414; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_415; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_416; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_417; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_418; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_419; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_420; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_421; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_422; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_423; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_424; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_425; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_426; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_427; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_428; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_429; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_430; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_431; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_432; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_433; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_434; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_435; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_436; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_437; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_438; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_439; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_440; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_441; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_442; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_443; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_444; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_445; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_446; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_447; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_448; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_449; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_450; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_451; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_452; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_453; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_454; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_455; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_456; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_457; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_458; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_459; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_460; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_461; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_462; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_463; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_464; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_465; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_466; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_467; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_468; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_469; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_470; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_471; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_472; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_473; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_474; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_475; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_476; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_477; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_478; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_479; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_480; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_481; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_482; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_483; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_484; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_485; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_486; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_487; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_488; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_489; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_490; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_491; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_492; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_493; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_494; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_495; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_496; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_497; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_498; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_499; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_500; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_501; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_502; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_503; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_504; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_505; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_506; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_507; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_508; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_509; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_510; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_511; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_512; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_513; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_514; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_515; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_516; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_517; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_518; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_519; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_520; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_521; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_522; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_523; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_524; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_525; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_526; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_527; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_528; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_529; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_530; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_531; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_532; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_533; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_534; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_535; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_536; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_537; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_538; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_539; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_540; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_541; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_542; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_543; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_544; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_545; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_546; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_547; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_548; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_549; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_550; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_551; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_552; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_553; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_554; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_555; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_556; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_557; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_558; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_559; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_560; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_561; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_562; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_563; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_564; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_565; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_566; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_567; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_568; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_569; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_570; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_571; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_572; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_573; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_574; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_575; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_576; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_577; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_578; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_579; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_580; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_581; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_582; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_583; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_584; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_585; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_586; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_587; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_588; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_589; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_590; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_591; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_592; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_593; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_594; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_595; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_596; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_597; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_598; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_599; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_600; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_601; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_602; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_603; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_604; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_605; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_606; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_607; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_608; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_609; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_610; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_611; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_612; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_613; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_614; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_615; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_616; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_617; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_618; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_619; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_620; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_621; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_622; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_623; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_624; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_625; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_626; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_627; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_628; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_629; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_630; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_631; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_632; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_633; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_634; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_635; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_636; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_637; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_638; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_639; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_640; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_641; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_642; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_643; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_644; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_645; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_646; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_647; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_648; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_649; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_650; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_651; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_652; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_653; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_654; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_655; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_656; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_657; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_658; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_659; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_660; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_661; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_662; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_663; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_664; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_665; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_666; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_667; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_668; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_669; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_670; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_671; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_672; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_673; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_674; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_675; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_676; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_677; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_678; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_679; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_680; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_681; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_682; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_683; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_684; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_685; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_686; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_687; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_688; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_689; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_690; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_691; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_692; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_693; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_694; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_695; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_696; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_697; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_698; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_699; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_700; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_701; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_702; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_703; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_704; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_705; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_706; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_707; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_708; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_709; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_710; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_711; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_712; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_713; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_714; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_715; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_716; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_717; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_718; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_719; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_720; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_721; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_722; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_723; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_724; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_725; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_726; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_727; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_728; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_729; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_730; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_731; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_732; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_733; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_734; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_735; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_736; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_737; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_738; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_739; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_740; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_741; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_742; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_743; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_744; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_745; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_746; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_747; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_748; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_749; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_750; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_751; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_752; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_753; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_754; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_755; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_756; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_757; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_758; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_759; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_760; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_761; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_762; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_763; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_764; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_765; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_766; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_767; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_768; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_769; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_770; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_771; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_772; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_773; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_774; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_775; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_776; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_777; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_778; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_779; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_780; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_781; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_782; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_783; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_784; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_785; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_786; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_787; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_788; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_789; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_790; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_791; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_792; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_793; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_794; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_795; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_796; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_797; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_798; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_799; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_800; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_801; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_802; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_803; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_804; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_805; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_806; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_807; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_808; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_809; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_810; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_811; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_812; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_813; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_814; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_815; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_816; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_817; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_818; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_819; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_820; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_821; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_822; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_823; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_824; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_825; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_826; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_827; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_828; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_829; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_830; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_831; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_832; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_833; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_834; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_835; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_836; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_837; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_838; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_839; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_840; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_841; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_842; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_843; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_844; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_845; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_846; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_847; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_848; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_849; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_850; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_851; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_852; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_853; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_854; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_855; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_856; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_857; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_858; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_859; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_860; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_861; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_862; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_863; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_864; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_865; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_866; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_867; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_868; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_869; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_870; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_871; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_872; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_873; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_874; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_875; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_876; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_877; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_878; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_879; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_880; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_881; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_882; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_883; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_884; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_885; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_886; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_887; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_888; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_889; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_890; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_891; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_892; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_893; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_894; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_895; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_896; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_897; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_898; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_899; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_900; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_901; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_902; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_903; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_904; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_905; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_906; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_907; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_908; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_909; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_910; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_911; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_912; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_913; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_914; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_915; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_916; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_917; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_918; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_919; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_920; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_921; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_922; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_923; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_924; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_925; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_926; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_927; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_928; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_929; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_930; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_931; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_932; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_933; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_934; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_935; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_936; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_937; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_938; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_939; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_940; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_941; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_942; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_943; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_944; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_945; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_946; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_947; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_948; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_949; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_950; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_951; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_952; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_953; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_954; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_955; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_956; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_957; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_958; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_959; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_960; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_961; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_962; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_963; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_964; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_965; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_966; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_967; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_968; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_969; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_970; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_971; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_972; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_973; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_974; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_975; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_976; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_977; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_978; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_979; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_980; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_981; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_982; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_983; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_984; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_985; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_986; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_987; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_988; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_989; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_990; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_991; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_992; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_993; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_994; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_995; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_996; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_997; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_998; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_999; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1000; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1001; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1002; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1003; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1004; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1005; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1006; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1007; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1008; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1009; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1010; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1011; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1012; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1013; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1014; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1015; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1016; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1017; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1018; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1019; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1020; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1021; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1022; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1023; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1024; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1025; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1026; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1027; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1028; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1029; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1030; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1031; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1032; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1033; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1034; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1035; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1036; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1037; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1038; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1039; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1040; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1041; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1042; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1043; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1044; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1045; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1046; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1047; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1048; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1049; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1050; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1051; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1052; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1053; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1054; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1055; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1056; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1057; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1058; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1059; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1060; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1061; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1062; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1063; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1064; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1065; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1066; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1067; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1068; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1069; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1070; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1071; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1072; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1073; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1074; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1075; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1076; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1077; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1078; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1079; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1080; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1081; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1082; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1083; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1084; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1085; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1086; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1087; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1088; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1089; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1090; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1091; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1092; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1093; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1094; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1095; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1096; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1097; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1098; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1099; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1100; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1101; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1102; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1103; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1104; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1105; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1106; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1107; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1108; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1109; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1110; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1111; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1112; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1113; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1114; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1115; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1116; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1117; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1118; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1119; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1120; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1121; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1122; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1123; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1124; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1125; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1126; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1127; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1128; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1129; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1130; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1131; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1132; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1133; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1134; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1135; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1136; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1137; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1138; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1139; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1140; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1141; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1142; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1143; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1144; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1145; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1146; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1147; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1148; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1149; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1150; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1151; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1152; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1153; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1154; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1155; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1156; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1157; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1158; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1159; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1160; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1161; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1162; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1163; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1164; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1165; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1166; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1167; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1168; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1169; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1170; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1171; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1172; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1173; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1174; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1175; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1176; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1177; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1178; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1179; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1180; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1181; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1182; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1183; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1184; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1185; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1186; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1187; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1188; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1189; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1190; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1191; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1192; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1193; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1194; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1195; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1196; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1197; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1198; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1199; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1200; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1201; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1202; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1203; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1204; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1205; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1206; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1207; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1208; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1209; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1210; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1211; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1212; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1213; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1214; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1215; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1216; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1217; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1218; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1219; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1220; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1221; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1222; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1223; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1224; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1225; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1226; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1227; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1228; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1229; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1230; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1231; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1232; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1233; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1234; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1235; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1236; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1237; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1238; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1239; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1240; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1241; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1242; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1243; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1244; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1245; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1246; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1247; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1248; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1249; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1250; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1251; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1252; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1253; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1254; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1255; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1256; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1257; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1258; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1259; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1260; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1261; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1262; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1263; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1264; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1265; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1266; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1267; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1268; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1269; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1270; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1271; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1272; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1273; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1274; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1275; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1276; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1277; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1278; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1279; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1280; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1281; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1282; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1283; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1284; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1285; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1286; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1287; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1288; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1289; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1290; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1291; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1292; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1293; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1294; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1295; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1296; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1297; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1298; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1299; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1300; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1301; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1302; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1303; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1304; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1305; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1306; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1307; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1308; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1309; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1310; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1311; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1312; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1313; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1314; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1315; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1316; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1317; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1318; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1319; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1320; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1321; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1322; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1323; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1324; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1325; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1326; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1327; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1328; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1329; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1330; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1331; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1332; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1333; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1334; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1335; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1336; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1337; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1338; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1339; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1340; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1341; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1342; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1343; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1344; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1345; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1346; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1347; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1348; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1349; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1350; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1351; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1352; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1353; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1354; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1355; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1356; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1357; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1358; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1359; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1360; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1361; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1362; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1363; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1364; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1365; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1366; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1367; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1368; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1369; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1370; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1371; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1372; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1373; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1374; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1375; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1376; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1377; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1378; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1379; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1380; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1381; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1382; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1383; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1384; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1385; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1386; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1387; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1388; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1389; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1390; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1391; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1392; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1393; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1394; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1395; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1396; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1397; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1398; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1399; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1400; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1401; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1402; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1403; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1404; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1405; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1406; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1407; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1408; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1409; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1410; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1411; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1412; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1413; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1414; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1415; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1416; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1417; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1418; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1419; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1420; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1421; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1422; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1423; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1424; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1425; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1426; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1427; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1428; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1429; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1430; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1431; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1432; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1433; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1434; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1435; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1436; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1437; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1438; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1439; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1440; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1441; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1442; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1443; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1444; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1445; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1446; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1447; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1448; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1449; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1450; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1451; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1452; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1453; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1454; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1455; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1456; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1457; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1458; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1459; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1460; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1461; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1462; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1463; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1464; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1465; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1466; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1467; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1468; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1469; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1470; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1471; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1472; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1473; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1474; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1475; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1476; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1477; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1478; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1479; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1480; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1481; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1482; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1483; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1484; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1485; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1486; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1487; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1488; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1489; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1490; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1491; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1492; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1493; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1494; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1495; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1496; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1497; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1498; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1499; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1500; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1501; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1502; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1503; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1504; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1505; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1506; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1507; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1508; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1509; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1510; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1511; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1512; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1513; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1514; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1515; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1516; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1517; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1518; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1519; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1520; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1521; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1522; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1523; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1524; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1525; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1526; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1527; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1528; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1529; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1530; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1531; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1532; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1533; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1534; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1535; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1536; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1537; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1538; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1539; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1540; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1541; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1542; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1543; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1544; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1545; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1546; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1547; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1548; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1549; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1550; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1551; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1552; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1553; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1554; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1555; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1556; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1557; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1558; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1559; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1560; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1561; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1562; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1563; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1564; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1565; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1566; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1567; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1568; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1569; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1570; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1571; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1572; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1573; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1574; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1575; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1576; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1577; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1578; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1579; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1580; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1581; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1582; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1583; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1584; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1585; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1586; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1587; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1588; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1589; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1590; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1591; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1592; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1593; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1594; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1595; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1596; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1597; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1598; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1599; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1600; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1601; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1602; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1603; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1604; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1605; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1606; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1607; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1608; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1609; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1610; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1611; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1612; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1613; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1614; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1615; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1616; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1617; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1618; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1619; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1620; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1621; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1622; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1623; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1624; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1625; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1626; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1627; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1628; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1629; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1630; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1631; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1632; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1633; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1634; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1635; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1636; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1637; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1638; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1639; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1640; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1641; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1642; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1643; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1644; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1645; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1646; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1647; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1648; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1649; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1650; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1651; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1652; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1653; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1654; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1655; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1656; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1657; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1658; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1659; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1660; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1661; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1662; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1663; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1664; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1665; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1666; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1667; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1668; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1669; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1670; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1671; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1672; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1673; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1674; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1675; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1676; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1677; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1678; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1679; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1680; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1681; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1682; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1683; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1684; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1685; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1686; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1687; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1688; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1689; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1690; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1691; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1692; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1693; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1694; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1695; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1696; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1697; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1698; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1699; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1700; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1701; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1702; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1703; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1704; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1705; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1706; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1707; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1708; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1709; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1710; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1711; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1712; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1713; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1714; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1715; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1716; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1717; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1718; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1719; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1720; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1721; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1722; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1723; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1724; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1725; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1726; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1727; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1728; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1729; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1730; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1731; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1732; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1733; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1734; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1735; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1736; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1737; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1738; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1739; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1740; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1741; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1742; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1743; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1744; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1745; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1746; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1747; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1748; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1749; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1750; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1751; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1752; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1753; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1754; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1755; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1756; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1757; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1758; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1759; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1760; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1761; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1762; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1763; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1764; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1765; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1766; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1767; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1768; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1769; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1770; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1771; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1772; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1773; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1774; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1775; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1776; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1777; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1778; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1779; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1780; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1781; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1782; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1783; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1784; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1785; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1786; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1787; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1788; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1789; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1790; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1791; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1792; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1793; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1794; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1795; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1796; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1797; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1798; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1799; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1800; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1801; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1802; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1803; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1804; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1805; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1806; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1807; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1808; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1809; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1810; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1811; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1812; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1813; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1814; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1815; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1816; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1817; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1818; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1819; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1820; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1821; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1822; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1823; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1824; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1825; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1826; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1827; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1828; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1829; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1830; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1831; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1832; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1833; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1834; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1835; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1836; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1837; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1838; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1839; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1840; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1841; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1842; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1843; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1844; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1845; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1846; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1847; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1848; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1849; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1850; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1851; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1852; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1853; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1854; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1855; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1856; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1857; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1858; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1859; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1860; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1861; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1862; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1863; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1864; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1865; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1866; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1867; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1868; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1869; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1870; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1871; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1872; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1873; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1874; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1875; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1876; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1877; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1878; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1879; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1880; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1881; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1882; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1883; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1884; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1885; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1886; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1887; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1888; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1889; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1890; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1891; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1892; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1893; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1894; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1895; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1896; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1897; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1898; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1899; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1900; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1901; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1902; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1903; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1904; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1905; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1906; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1907; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1908; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1909; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1910; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1911; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1912; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1913; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1914; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1915; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1916; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1917; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1918; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1919; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1920; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1921; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1922; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1923; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1924; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1925; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1926; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1927; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1928; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1929; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1930; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1931; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1932; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1933; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1934; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1935; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1936; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1937; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1938; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1939; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1940; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1941; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1942; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1943; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1944; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1945; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1946; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1947; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1948; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1949; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1950; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1951; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1952; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1953; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1954; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1955; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1956; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1957; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1958; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1959; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1960; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1961; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1962; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1963; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1964; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1965; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1966; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1967; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1968; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1969; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1970; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1971; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1972; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1973; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1974; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1975; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1976; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1977; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1978; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1979; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1980; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1981; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1982; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1983; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1984; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1985; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1986; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1987; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1988; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1989; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1990; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1991; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1992; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1993; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1994; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1995; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1996; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1997; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1998; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_1999; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2000; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2001; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2002; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2003; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2004; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2005; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2006; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2007; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2008; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2009; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2010; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2011; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2012; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2013; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2014; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2015; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2016; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2017; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2018; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2019; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2020; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2021; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2022; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2023; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2024; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2025; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2026; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2027; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2028; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2029; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2030; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2031; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2032; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2033; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2034; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2035; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2036; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2037; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2038; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2039; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2040; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2041; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2042; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2043; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2044; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2045; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2046; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2047; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2048; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2049; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2050; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2051; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2052; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2053; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2054; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2055; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2056; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2057; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2058; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2059; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2060; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2061; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2062; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2063; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2064; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2065; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2066; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2067; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2068; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2069; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2070; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2071; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2072; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2073; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2074; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2075; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2076; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2077; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2078; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2079; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2080; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2081; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2082; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2083; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2084; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2085; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2086; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2087; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2088; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2089; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2090; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2091; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2092; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2093; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2094; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2095; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2096; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2097; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2098; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2099; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2100; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2101; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2102; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2103; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2104; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2105; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2106; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2107; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2108; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2109; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2110; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2111; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2112; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2113; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2114; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2115; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2116; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2117; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2118; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2119; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2120; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2121; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2122; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2123; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2124; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2125; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire  _GEN_2126; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  wire [3:0] _GEN_4175; // @[TLSimpleL2.scala 326:40:freechips.rocketchip.system.DefaultConfig.fir@223412.4]
  wire [15:0] _T_604_0; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221284.4]
  wire [15:0] _T_604_1; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221285.4]
  wire [15:0] _T_604_2; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221286.4]
  wire [15:0] _T_604_3; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221287.4]
  wire [15:0] _T_604_4; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221288.4]
  wire [15:0] _T_604_5; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221289.4]
  wire [15:0] _T_604_6; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221290.4]
  wire [15:0] _T_604_7; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221291.4]
  wire [15:0] _T_604_8; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221292.4]
  wire [15:0] _T_604_9; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221293.4]
  wire [15:0] _T_604_10; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221294.4]
  wire [15:0] _T_604_11; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221295.4]
  wire [15:0] _T_604_12; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221296.4]
  wire [15:0] _T_604_13; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221297.4]
  wire [15:0] _T_604_14; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221298.4]
  wire [15:0] _T_604_15; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221299.4]
  wire [3:0] _T_663_0; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221335.4]
  wire [3:0] _T_663_1; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221336.4]
  wire [3:0] _T_663_2; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221337.4]
  wire [3:0] _T_663_3; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221338.4]
  wire [3:0] _T_663_4; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221339.4]
  wire [3:0] _T_663_5; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221340.4]
  wire [3:0] _T_663_6; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221341.4]
  wire [3:0] _T_663_7; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221342.4]
  wire [3:0] _T_663_8; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221343.4]
  wire [3:0] _T_663_9; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221344.4]
  wire [3:0] _T_663_10; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221345.4]
  wire [3:0] _T_663_11; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221346.4]
  wire [3:0] _T_663_12; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221347.4]
  wire [3:0] _T_663_13; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221348.4]
  wire [3:0] _T_663_14; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221349.4]
  wire [3:0] _T_663_15; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221350.4]
  wire [15:0] _T_13044; // @[TLSimpleL2.scala 337:21:freechips.rocketchip.system.DefaultConfig.fir@223422.4]
  wire  _T_13045; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223423.4]
  wire  _T_13046; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223424.4]
  wire  _T_13047; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223425.4]
  wire  _T_13048; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223426.4]
  wire  _T_13049; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223427.4]
  wire  _T_13050; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223428.4]
  wire  _T_13051; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223429.4]
  wire  _T_13052; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223430.4]
  wire  _T_13053; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223431.4]
  wire  _T_13054; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223432.4]
  wire  _T_13055; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223433.4]
  wire  _T_13056; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223434.4]
  wire  _T_13057; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223435.4]
  wire  _T_13058; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223436.4]
  wire  _T_13059; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223437.4]
  wire  _T_13060; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223438.4]
  wire  _T_13083; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223457.4]
  wire  _T_13084; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223458.4]
  wire  _T_13085; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223459.4]
  wire  _T_13086; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223460.4]
  wire  _T_13087; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223461.4]
  wire  _T_13088; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223462.4]
  wire  _T_13089; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223463.4]
  wire  _T_13090; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223464.4]
  wire  _T_13091; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223465.4]
  wire  _T_13092; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223466.4]
  wire  _T_13093; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223467.4]
  wire  _T_13094; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223468.4]
  wire  _T_13095; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223469.4]
  wire  _T_13096; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223470.4]
  wire  _T_13097; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223471.4]
  wire  _T_13098; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223472.4]
  wire  _T_13099; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223473.4]
  wire  _T_13100; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223474.4]
  wire  _T_13101; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223475.4]
  wire  _T_13102; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223476.4]
  wire  _T_13103; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223477.4]
  wire  _T_13104; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223478.4]
  wire  _T_13105; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223479.4]
  wire  _T_13106; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223480.4]
  wire  _T_13107; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223481.4]
  wire  _T_13108; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223482.4]
  wire  _T_13109; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223483.4]
  wire  _T_13110; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223484.4]
  wire  _T_13111; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223485.4]
  wire  _T_13112; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223486.4]
  wire  _T_13113; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223487.4]
  wire  _T_13114; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223488.4]
  wire [1:0] _T_13137; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223507.4]
  wire [1:0] _T_13138; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223508.4]
  wire [3:0] _T_13139; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223509.4]
  wire [1:0] _T_13140; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223510.4]
  wire [1:0] _T_13141; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223511.4]
  wire [3:0] _T_13142; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223512.4]
  wire [7:0] _T_13143; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223513.4]
  wire [1:0] _T_13144; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223514.4]
  wire [1:0] _T_13145; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223515.4]
  wire [3:0] _T_13146; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223516.4]
  wire [1:0] _T_13147; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223517.4]
  wire [1:0] _T_13148; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223518.4]
  wire [3:0] _T_13149; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223519.4]
  wire [7:0] _T_13150; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223520.4]
  wire [15:0] _T_13151; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223521.4]
  wire  _T_13152; // @[TLSimpleL2.scala 340:31:freechips.rocketchip.system.DefaultConfig.fir@223522.4]
  wire  _T_13153; // @[TLSimpleL2.scala 341:26:freechips.rocketchip.system.DefaultConfig.fir@223523.4]
  wire  _T_13154; // @[TLSimpleL2.scala 342:27:freechips.rocketchip.system.DefaultConfig.fir@223524.4]
  wire  _T_13155; // @[TLSimpleL2.scala 343:23:freechips.rocketchip.system.DefaultConfig.fir@223525.4]
  wire  _T_13156; // @[TLSimpleL2.scala 343:28:freechips.rocketchip.system.DefaultConfig.fir@223526.4]
  wire  _T_13158; // @[TLSimpleL2.scala 344:29:freechips.rocketchip.system.DefaultConfig.fir@223528.4]
  wire  _T_13162; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223536.4]
  wire  _T_13163; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223540.4]
  wire [1:0] _GEN_6261; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223541.4]
  wire  _T_13164; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223544.4]
  wire [1:0] _GEN_6262; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223545.4]
  wire  _T_13165; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223548.4]
  wire [2:0] _GEN_6263; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223549.4]
  wire  _T_13166; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223552.4]
  wire [2:0] _GEN_6264; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223553.4]
  wire  _T_13167; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223556.4]
  wire [2:0] _GEN_6265; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223557.4]
  wire  _T_13168; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223560.4]
  wire [2:0] _GEN_6266; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223561.4]
  wire  _T_13169; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223564.4]
  wire [3:0] _GEN_6267; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223565.4]
  wire  _T_13170; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223568.4]
  wire [3:0] _GEN_6268; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223569.4]
  wire  _T_13171; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223572.4]
  wire [3:0] _GEN_6269; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223573.4]
  wire  _T_13172; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223576.4]
  wire [3:0] _GEN_6270; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223577.4]
  wire  _T_13173; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223580.4]
  wire [3:0] _GEN_6271; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223581.4]
  wire  _T_13174; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223584.4]
  wire [3:0] _GEN_6272; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223585.4]
  wire  _T_13175; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223588.4]
  wire [3:0] _GEN_6273; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223589.4]
  wire  _T_13176; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223592.4]
  wire [3:0] _GEN_6274; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223593.4]
  wire [15:0] _T_13177; // @[TLSimpleL2.scala 351:42:freechips.rocketchip.system.DefaultConfig.fir@223597.4]
  wire  _T_13178; // @[TLSimpleL2.scala 351:55:freechips.rocketchip.system.DefaultConfig.fir@223598.4]
  wire  _T_13180; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223600.4]
  wire  _T_13181; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223601.4]
  wire  _T_13182; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223602.4]
  wire  _T_13183; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223603.4]
  wire  _T_13184; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223604.4]
  wire  _T_13185; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223605.4]
  wire  _T_13186; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223606.4]
  wire  _T_13187; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223607.4]
  wire  _T_13188; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223608.4]
  wire  _T_13189; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223609.4]
  wire  _T_13190; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223610.4]
  wire  _T_13191; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223611.4]
  wire  _T_13192; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223612.4]
  wire  _T_13193; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223613.4]
  wire  _T_13194; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223614.4]
  wire [3:0] _T_13196; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223616.4]
  wire [3:0] _T_13197; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223617.4]
  wire [3:0] _T_13198; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223618.4]
  wire [3:0] _T_13199; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223619.4]
  wire [3:0] _T_13200; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223620.4]
  wire [3:0] _T_13201; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223621.4]
  wire [3:0] _T_13202; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223622.4]
  wire [3:0] _T_13203; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223623.4]
  wire [3:0] _T_13204; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223624.4]
  wire [3:0] _T_13205; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223625.4]
  wire [3:0] _T_13206; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223626.4]
  wire [3:0] _T_13207; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223627.4]
  wire [3:0] _T_13208; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223628.4]
  wire [3:0] _T_13209; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223629.4]
  wire [3:0] _T_13210; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223630.4]
  wire  _T_13211; // @[TLSimpleL2.scala 352:23:freechips.rocketchip.system.DefaultConfig.fir@223631.4]
  wire  _T_13212; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223632.4]
  wire  _T_13213; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223633.4]
  wire  _T_13214; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223634.4]
  wire  _T_13215; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223635.4]
  wire  _T_13216; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223636.4]
  wire  _T_13217; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223637.4]
  wire  _T_13218; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223638.4]
  wire  _T_13219; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223639.4]
  wire  _T_13220; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223640.4]
  wire  _T_13221; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223641.4]
  wire  _T_13222; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223642.4]
  wire  _T_13223; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223643.4]
  wire  _T_13224; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223644.4]
  wire  _T_13225; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223645.4]
  wire  _T_13226; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223646.4]
  wire [3:0] _T_13228; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223648.4]
  wire [3:0] _T_13229; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223649.4]
  wire [3:0] _T_13230; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223650.4]
  wire [3:0] _T_13231; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223651.4]
  wire [3:0] _T_13232; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223652.4]
  wire [3:0] _T_13233; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223653.4]
  wire [3:0] _T_13234; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223654.4]
  wire [3:0] _T_13235; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223655.4]
  wire [3:0] _T_13236; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223656.4]
  wire [3:0] _T_13237; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223657.4]
  wire [3:0] _T_13238; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223658.4]
  wire [3:0] _T_13239; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223659.4]
  wire [3:0] _T_13240; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223660.4]
  wire [3:0] _T_13241; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223661.4]
  wire [3:0] _T_13242; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223662.4]
  wire [3:0] _T_13243; // @[TLSimpleL2.scala 352:12:freechips.rocketchip.system.DefaultConfig.fir@223663.4]
  wire [3:0] _T_13244; // @[TLSimpleL2.scala 351:25:freechips.rocketchip.system.DefaultConfig.fir@223664.4]
  reg [14:0] _T_13304_0; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2111;
  reg [14:0] _T_13304_1; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2112;
  reg [14:0] _T_13304_2; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2113;
  reg [14:0] _T_13304_3; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2114;
  reg [14:0] _T_13304_4; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2115;
  reg [14:0] _T_13304_5; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2116;
  reg [14:0] _T_13304_6; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2117;
  reg [14:0] _T_13304_7; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2118;
  reg [14:0] _T_13304_8; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2119;
  reg [14:0] _T_13304_9; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2120;
  reg [14:0] _T_13304_10; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2121;
  reg [14:0] _T_13304_11; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2122;
  reg [14:0] _T_13304_12; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2123;
  reg [14:0] _T_13304_13; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2124;
  reg [14:0] _T_13304_14; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2125;
  reg [14:0] _T_13304_15; // @[TLSimpleL2.scala 354:34:freechips.rocketchip.system.DefaultConfig.fir@223683.4]
  reg [31:0] _RAND_2126;
  wire [14:0] _GEN_6276; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6277; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6278; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6279; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6280; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6281; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6282; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6283; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6284; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6285; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6286; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6287; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6288; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [14:0] _GEN_6289; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  wire [15:0] _T_13367; // @[TLSimpleL2.scala 365:40:freechips.rocketchip.system.DefaultConfig.fir@223688.4]
  wire  _T_13368; // @[TLSimpleL2.scala 365:40:freechips.rocketchip.system.DefaultConfig.fir@223689.4]
  wire [15:0] _T_13369; // @[TLSimpleL2.scala 365:66:freechips.rocketchip.system.DefaultConfig.fir@223690.4]
  wire  _T_13370; // @[TLSimpleL2.scala 365:66:freechips.rocketchip.system.DefaultConfig.fir@223691.4]
  wire  _T_13371; // @[TLSimpleL2.scala 365:51:freechips.rocketchip.system.DefaultConfig.fir@223692.4]
  wire [16:0] _T_13373; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223693.4]
  wire [15:0] _GEN_6292; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6293; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6294; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6295; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6296; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6297; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6298; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6299; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6300; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6301; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6302; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6303; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6304; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6305; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [15:0] _GEN_6306; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire [32:0] _T_13374; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  wire  _T_13375; // @[TLSimpleL2.scala 369:43:freechips.rocketchip.system.DefaultConfig.fir@223695.4]
  wire  _T_13376; // @[TLSimpleL2.scala 370:49:freechips.rocketchip.system.DefaultConfig.fir@223696.4]
  wire  _T_13377; // @[TLSimpleL2.scala 370:46:freechips.rocketchip.system.DefaultConfig.fir@223697.4]
  wire  _T_13378; // @[TLSimpleL2.scala 371:45:freechips.rocketchip.system.DefaultConfig.fir@223698.4]
  wire  _T_13380; // @[TLSimpleL2.scala 372:48:freechips.rocketchip.system.DefaultConfig.fir@223700.4]
  wire  _T_13381; // @[TLSimpleL2.scala 374:37:freechips.rocketchip.system.DefaultConfig.fir@223701.4]
  wire  _T_13382; // @[TLSimpleL2.scala 374:50:freechips.rocketchip.system.DefaultConfig.fir@223702.4]
  wire  _T_13383; // @[TLSimpleL2.scala 374:73:freechips.rocketchip.system.DefaultConfig.fir@223703.4]
  wire  _T_13385; // @[TLSimpleL2.scala 395:31:freechips.rocketchip.system.DefaultConfig.fir@223717.6]
  wire  _T_13387; // @[TLSimpleL2.scala 395:15:freechips.rocketchip.system.DefaultConfig.fir@223719.6]
  wire  _T_13388; // @[TLSimpleL2.scala 395:15:freechips.rocketchip.system.DefaultConfig.fir@223720.6]
  wire  _T_13392; // @[TLSimpleL2.scala 399:45:freechips.rocketchip.system.DefaultConfig.fir@223732.8]
  wire [3:0] _GEN_6307; // @[TLSimpleL2.scala 399:73:freechips.rocketchip.system.DefaultConfig.fir@223733.8]
  wire [3:0] _GEN_6308; // @[TLSimpleL2.scala 397:85:freechips.rocketchip.system.DefaultConfig.fir@223728.6]
  wire [3:0] _GEN_6309; // @[TLSimpleL2.scala 376:35:freechips.rocketchip.system.DefaultConfig.fir@223705.4]
  wire [3:0] _T_13418; // @[TLSimpleL2.scala 419:27:freechips.rocketchip.system.DefaultConfig.fir@223812.4]
  wire  _T_13424; // @[TLSimpleL2.scala 422:15:freechips.rocketchip.system.DefaultConfig.fir@223819.6]
  wire [15:0] _T_13425; // @[TLSimpleL2.scala 423:40:freechips.rocketchip.system.DefaultConfig.fir@223821.8]
  wire [15:0] _T_13426; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223825.8]
  wire [15:0] _T_13428; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223827.8]
  wire [15:0] _T_13429; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223828.8]
  wire [15:0] _T_13430; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223829.8]
  wire [15:0] _GEN_6310; // @[TLSimpleL2.scala 422:50:freechips.rocketchip.system.DefaultConfig.fir@223820.6]
  wire  _T_13454; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223836.4]
  wire [15:0] _T_13455; // @[TLSimpleL2.scala 437:55:freechips.rocketchip.system.DefaultConfig.fir@223839.6]
  wire  _T_13456; // @[TLSimpleL2.scala 437:55:freechips.rocketchip.system.DefaultConfig.fir@223840.6]
  wire  _T_13457; // @[TLSimpleL2.scala 438:16:freechips.rocketchip.system.DefaultConfig.fir@223841.6]
  wire  _T_13458; // @[TLSimpleL2.scala 437:32:freechips.rocketchip.system.DefaultConfig.fir@223842.6]
  wire  _T_13460; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223850.6]
  wire  _GEN_6312; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  wire  _GEN_6313; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  wire [15:0] _GEN_6314; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  wire [3:0] _GEN_6315; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  wire  _T_13461; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223855.4]
  wire  _T_13462; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223857.4]
  wire  _T_13468; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223871.6]
  wire  _GEN_6316; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  wire  _GEN_6317; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  wire [15:0] _GEN_6318; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  wire [3:0] _GEN_6319; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  wire  _T_13469; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223876.4]
  wire  _T_13470; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223878.4]
  wire  _T_13476; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223892.6]
  wire  _GEN_6320; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  wire  _GEN_6321; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  wire [15:0] _GEN_6322; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  wire [3:0] _GEN_6323; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  wire  _T_13477; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223897.4]
  wire  _T_13478; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223899.4]
  wire  _T_13484; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223913.6]
  wire  _GEN_6324; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  wire  _GEN_6325; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  wire [15:0] _GEN_6326; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  wire [3:0] _GEN_6327; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  wire  _T_13485; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223918.4]
  wire  _T_13486; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223920.4]
  wire  _T_13492; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223934.6]
  wire  _GEN_6328; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  wire  _GEN_6329; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  wire [15:0] _GEN_6330; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  wire [3:0] _GEN_6331; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  wire  _T_13493; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223939.4]
  wire  _T_13494; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223941.4]
  wire  _T_13500; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223955.6]
  wire  _GEN_6332; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  wire  _GEN_6333; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  wire [15:0] _GEN_6334; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  wire [3:0] _GEN_6335; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  wire  _T_13501; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223960.4]
  wire  _T_13502; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223962.4]
  wire  _T_13508; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223976.6]
  wire  _GEN_6336; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  wire  _GEN_6337; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  wire [15:0] _GEN_6338; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  wire [3:0] _GEN_6339; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  wire  _T_13509; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223981.4]
  wire  _T_13510; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223983.4]
  wire  _T_13516; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223997.6]
  wire  _GEN_6340; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  wire  _GEN_6341; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  wire [15:0] _GEN_6342; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  wire [3:0] _GEN_6343; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  wire  _T_13517; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224002.4]
  wire  _T_13518; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224004.4]
  wire  _T_13524; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224018.6]
  wire  _GEN_6344; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  wire  _GEN_6345; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  wire [15:0] _GEN_6346; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  wire [3:0] _GEN_6347; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  wire  _T_13525; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224023.4]
  wire  _T_13526; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224025.4]
  wire  _T_13532; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224039.6]
  wire  _GEN_6348; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  wire  _GEN_6349; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  wire [15:0] _GEN_6350; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  wire [3:0] _GEN_6351; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  wire  _T_13533; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224044.4]
  wire  _T_13534; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224046.4]
  wire  _T_13540; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224060.6]
  wire  _GEN_6352; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  wire  _GEN_6353; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  wire [15:0] _GEN_6354; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  wire [3:0] _GEN_6355; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  wire  _T_13541; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224065.4]
  wire  _T_13542; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224067.4]
  wire  _T_13548; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224081.6]
  wire  _GEN_6356; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  wire  _GEN_6357; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  wire [15:0] _GEN_6358; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  wire [3:0] _GEN_6359; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  wire  _T_13549; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224086.4]
  wire  _T_13550; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224088.4]
  wire  _T_13556; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224102.6]
  wire  _GEN_6360; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  wire  _GEN_6361; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  wire [15:0] _GEN_6362; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  wire [3:0] _GEN_6363; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  wire  _T_13557; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224107.4]
  wire  _T_13558; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224109.4]
  wire  _T_13564; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224123.6]
  wire  _GEN_6364; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  wire  _GEN_6365; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  wire [15:0] _GEN_6366; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  wire [3:0] _GEN_6367; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  wire  _T_13565; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224128.4]
  wire  _T_13566; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224130.4]
  wire  _T_13572; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224144.6]
  wire  _GEN_6368; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  wire  _GEN_6369; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  wire [15:0] _GEN_6370; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  wire [3:0] _GEN_6371; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  wire  _T_13573; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224149.4]
  wire  _T_13574; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224151.4]
  wire  _T_13580; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224165.6]
  wire  _GEN_6372; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  wire  _GEN_6373; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  wire [15:0] _GEN_6374; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  wire [3:0] _GEN_6375; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  wire  _T_13581; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224170.4]
  wire [12:0] _T_13583; // @[TLSimpleL2.scala 455:32:freechips.rocketchip.system.DefaultConfig.fir@224175.4]
  wire [15:0] _T_13435_0_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223845.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223853.6]
  wire [15:0] _T_13584_0_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_1_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223866.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223874.6]
  wire [15:0] _T_13584_1_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_2_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223887.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223895.6]
  wire [15:0] _T_13584_2_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_3_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223908.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223916.6]
  wire [15:0] _T_13584_3_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_4_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223929.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223937.6]
  wire [15:0] _T_13584_4_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_5_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223950.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223958.6]
  wire [15:0] _T_13584_5_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_6_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223971.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223979.6]
  wire [15:0] _T_13584_6_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_7_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223992.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224000.6]
  wire [15:0] _T_13584_7_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_8_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224013.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224021.6]
  wire [15:0] _T_13584_8_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_9_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224034.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224042.6]
  wire [15:0] _T_13584_9_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_10_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224055.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224063.6]
  wire [15:0] _T_13584_10_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_11_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224076.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224084.6]
  wire [15:0] _T_13584_11_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_12_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224097.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224105.6]
  wire [15:0] _T_13584_12_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_13_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224118.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224126.6]
  wire [15:0] _T_13584_13_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_14_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224139.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224147.6]
  wire [15:0] _T_13584_14_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [15:0] _T_13435_15_dsid; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224160.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224168.6]
  wire [15:0] _T_13584_15_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  wire [10:0] _T_13620; // @[:freechips.rocketchip.system.DefaultConfig.fir@224178.6]
  wire  _T_13659; // @[TLSimpleL2.scala 461:20:freechips.rocketchip.system.DefaultConfig.fir@224183.6]
  wire  _T_13660; // @[TLSimpleL2.scala 462:29:freechips.rocketchip.system.DefaultConfig.fir@224185.8]
  wire  _T_13662; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224187.8]
  wire  _T_13663; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224188.8]
  wire  _T_13666; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224195.8]
  wire  _T_13667; // @[TLSimpleL2.scala 465:38:freechips.rocketchip.system.DefaultConfig.fir@224196.8]
  wire [3:0] _GEN_6377; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6378; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6379; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6380; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6381; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6382; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6383; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6384; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6385; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6386; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6387; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6388; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6389; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6390; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire [3:0] _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire  _T_13668; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  wire  _T_13669; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224198.8]
  wire  _T_13670; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224199.8]
  wire [14:0] _GEN_6393; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6394; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6395; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6396; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6397; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6398; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6399; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6400; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6401; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6402; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6403; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6404; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6405; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6406; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _GEN_6407; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  wire [14:0] _T_13672; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224202.10]
  wire  _T_13673; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224206.10]
  wire  _T_13674; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224207.10]
  wire  _T_13675; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224208.10]
  wire  _T_13676; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224209.10]
  wire [14:0] _GEN_6409; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6410; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6411; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6412; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6413; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6414; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6415; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6416; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6417; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6418; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6419; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6420; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6421; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6422; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [14:0] _GEN_6423; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [15:0] _T_13677; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  wire [15:0] _T_13678; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224212.12]
  wire [14:0] _T_13679; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224213.12]
  wire  _T_13680; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224216.8]
  wire  _T_13682; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224218.8]
  wire  _T_13683; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224219.8]
  wire  _T_13684; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224220.8]
  wire  _T_13687; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224227.10]
  wire  _T_13688; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224228.10]
  wire  _T_13689; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224229.10]
  wire  _T_13690; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224230.10]
  wire  _T_13694; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224237.8]
  wire  _T_13696; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224239.8]
  wire  _T_13697; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224240.8]
  wire  _T_13698; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224241.8]
  wire  _T_13701; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224248.10]
  wire  _T_13702; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224249.10]
  wire  _T_13703; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224250.10]
  wire  _T_13704; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224251.10]
  wire  _T_13708; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224258.8]
  wire  _T_13710; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224260.8]
  wire  _T_13711; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224261.8]
  wire  _T_13712; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224262.8]
  wire  _T_13715; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224269.10]
  wire  _T_13716; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224270.10]
  wire  _T_13717; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224271.10]
  wire  _T_13718; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224272.10]
  wire  _T_13722; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224279.8]
  wire  _T_13724; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224281.8]
  wire  _T_13725; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224282.8]
  wire  _T_13726; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224283.8]
  wire  _T_13729; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224290.10]
  wire  _T_13730; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224291.10]
  wire  _T_13731; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224292.10]
  wire  _T_13732; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224293.10]
  wire  _T_13736; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224300.8]
  wire  _T_13738; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224302.8]
  wire  _T_13739; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224303.8]
  wire  _T_13740; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224304.8]
  wire  _T_13743; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224311.10]
  wire  _T_13744; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224312.10]
  wire  _T_13745; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224313.10]
  wire  _T_13746; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224314.10]
  wire  _T_13750; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224321.8]
  wire  _T_13752; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224323.8]
  wire  _T_13753; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224324.8]
  wire  _T_13754; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224325.8]
  wire  _T_13757; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224332.10]
  wire  _T_13758; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224333.10]
  wire  _T_13759; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224334.10]
  wire  _T_13760; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224335.10]
  wire  _T_13764; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224342.8]
  wire  _T_13766; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224344.8]
  wire  _T_13767; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224345.8]
  wire  _T_13768; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224346.8]
  wire  _T_13771; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224353.10]
  wire  _T_13772; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224354.10]
  wire  _T_13773; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224355.10]
  wire  _T_13774; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224356.10]
  wire  _T_13778; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224363.8]
  wire  _T_13780; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224365.8]
  wire  _T_13781; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224366.8]
  wire  _T_13782; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224367.8]
  wire  _T_13785; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224374.10]
  wire  _T_13786; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224375.10]
  wire  _T_13787; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224376.10]
  wire  _T_13788; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224377.10]
  wire  _T_13792; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224384.8]
  wire  _T_13794; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224386.8]
  wire  _T_13795; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224387.8]
  wire  _T_13796; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224388.8]
  wire  _T_13799; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224395.10]
  wire  _T_13800; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224396.10]
  wire  _T_13801; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224397.10]
  wire  _T_13802; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224398.10]
  wire  _T_13806; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224405.8]
  wire  _T_13808; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224407.8]
  wire  _T_13809; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224408.8]
  wire  _T_13810; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224409.8]
  wire  _T_13813; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224416.10]
  wire  _T_13814; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224417.10]
  wire  _T_13815; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224418.10]
  wire  _T_13816; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224419.10]
  wire  _T_13820; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224426.8]
  wire  _T_13822; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224428.8]
  wire  _T_13823; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224429.8]
  wire  _T_13824; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224430.8]
  wire  _T_13827; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224437.10]
  wire  _T_13828; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224438.10]
  wire  _T_13829; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224439.10]
  wire  _T_13830; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224440.10]
  wire  _T_13834; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224447.8]
  wire  _T_13836; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224449.8]
  wire  _T_13837; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224450.8]
  wire  _T_13838; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224451.8]
  wire  _T_13841; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224458.10]
  wire  _T_13842; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224459.10]
  wire  _T_13843; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224460.10]
  wire  _T_13844; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224461.10]
  wire  _T_13848; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224468.8]
  wire  _T_13850; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224470.8]
  wire  _T_13851; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224471.8]
  wire  _T_13852; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224472.8]
  wire  _T_13855; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224479.10]
  wire  _T_13856; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224480.10]
  wire  _T_13857; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224481.10]
  wire  _T_13858; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224482.10]
  wire  _T_13862; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224489.8]
  wire  _T_13864; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224491.8]
  wire  _T_13865; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224492.8]
  wire  _T_13866; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224493.8]
  wire  _T_13869; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224500.10]
  wire  _T_13870; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224501.10]
  wire  _T_13871; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224502.10]
  wire  _T_13872; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224503.10]
  wire  _T_13876; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224510.8]
  wire  _T_13878; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224512.8]
  wire  _T_13879; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224513.8]
  wire  _T_13880; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224514.8]
  wire  _T_13883; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224521.10]
  wire  _T_13884; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224522.10]
  wire  _T_13885; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224523.10]
  wire  _T_13886; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224524.10]
  wire [3:0] _T_13891; // @[TLSimpleL2.scala 481:30:freechips.rocketchip.system.DefaultConfig.fir@224536.4]
  reg [3:0] _T_13893; // @[TLSimpleL2.scala 483:34:freechips.rocketchip.system.DefaultConfig.fir@224537.4]
  reg [31:0] _RAND_2127;
  wire  _T_13895; // @[TLSimpleL2.scala 484:51:freechips.rocketchip.system.DefaultConfig.fir@224539.4]
  wire  _T_13896; // @[TLSimpleL2.scala 484:80:freechips.rocketchip.system.DefaultConfig.fir@224540.4]
  wire  _T_13897; // @[TLSimpleL2.scala 484:113:freechips.rocketchip.system.DefaultConfig.fir@224541.4]
  wire  _T_13898; // @[TLSimpleL2.scala 484:96:freechips.rocketchip.system.DefaultConfig.fir@224542.4]
  wire  _T_13899; // @[TLSimpleL2.scala 484:70:freechips.rocketchip.system.DefaultConfig.fir@224543.4]
  wire [13:0] _GEN_7028; // @[TLSimpleL2.scala 485:31:freechips.rocketchip.system.DefaultConfig.fir@224544.4]
  wire [13:0] _T_13900; // @[TLSimpleL2.scala 485:31:freechips.rocketchip.system.DefaultConfig.fir@224544.4]
  wire [13:0] _GEN_7029; // @[TLSimpleL2.scala 485:59:freechips.rocketchip.system.DefaultConfig.fir@224545.4]
  wire [13:0] _T_13901; // @[TLSimpleL2.scala 485:59:freechips.rocketchip.system.DefaultConfig.fir@224545.4]
  wire [3:0] _T_13909; // @[TLSimpleL2.scala 488:31:freechips.rocketchip.system.DefaultConfig.fir@224548.4]
  wire  _T_13912; // @[TLSimpleL2.scala 490:36:freechips.rocketchip.system.DefaultConfig.fir@224551.4]
  reg [2:0] value_1; // @[Counter.scala 26:33:freechips.rocketchip.system.DefaultConfig.fir@224757.4]
  reg [31:0] _RAND_2128;
  wire [13:0] _GEN_7031; // @[TLSimpleL2.scala 491:60:freechips.rocketchip.system.DefaultConfig.fir@224553.4]
  wire [13:0] _T_13914; // @[TLSimpleL2.scala 491:60:freechips.rocketchip.system.DefaultConfig.fir@224553.4]
  wire [3:0] _T_14156; // @[TLSimpleL2.scala 559:49:freechips.rocketchip.system.DefaultConfig.fir@224767.4]
  wire [2:0] _T_14157; // @[TLSimpleL2.scala 559:49:freechips.rocketchip.system.DefaultConfig.fir@224768.4]
  reg [63:0] _T_14075_7; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2129;
  reg [63:0] _T_14075_6; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2130;
  reg [63:0] _T_14075_5; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2131;
  reg [63:0] _T_14075_4; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2132;
  reg [63:0] _T_14075_3; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2133;
  reg [63:0] _T_14075_2; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2134;
  reg [63:0] _T_14075_1; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2135;
  reg [63:0] _T_14075_0; // @[TLSimpleL2.scala 515:25:freechips.rocketchip.system.DefaultConfig.fir@224666.4]
  reg [63:0] _RAND_2136;
  wire [63:0] _GEN_6968; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  wire [63:0] _GEN_6969; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  wire [63:0] _GEN_6970; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  wire [63:0] _GEN_6971; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  wire [63:0] _GEN_6972; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  wire [63:0] _GEN_6973; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  wire  _T_14020; // @[TLSimpleL2.scala 506:70:freechips.rocketchip.system.DefaultConfig.fir@224644.4]
  wire  _T_14021; // @[TLSimpleL2.scala 506:67:freechips.rocketchip.system.DefaultConfig.fir@224645.4]
  wire [63:0] _GEN_6883; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6884; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6885; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6886; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6887; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6888; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6889; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6890; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6891; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6892; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6893; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6894; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6895; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6896; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6897; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [63:0] _GEN_6898; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  wire [3:0] _T_14087; // @[TLSimpleL2.scala 517:40:freechips.rocketchip.system.DefaultConfig.fir@224669.6]
  wire [4:0] _T_14089; // @[TLSimpleL2.scala 521:36:freechips.rocketchip.system.DefaultConfig.fir@224674.6]
  wire [4:0] _T_14090; // @[TLSimpleL2.scala 521:36:freechips.rocketchip.system.DefaultConfig.fir@224675.6]
  wire [3:0] _T_14091; // @[TLSimpleL2.scala 521:36:freechips.rocketchip.system.DefaultConfig.fir@224676.6]
  wire [4:0] _T_14093; // @[TLSimpleL2.scala 521:57:freechips.rocketchip.system.DefaultConfig.fir@224678.6]
  wire [3:0] _T_14094; // @[TLSimpleL2.scala 521:57:freechips.rocketchip.system.DefaultConfig.fir@224679.6]
  wire [2:0] _T_14096; // @[:freechips.rocketchip.system.DefaultConfig.fir@224680.6]
  wire  _T_14097; // @[TLSimpleL2.scala 523:29:freechips.rocketchip.system.DefaultConfig.fir@224682.6]
  wire  _T_14098; // @[TLSimpleL2.scala 527:44:freechips.rocketchip.system.DefaultConfig.fir@224689.10]
  wire [3:0] _GEN_6908; // @[TLSimpleL2.scala 529:35:freechips.rocketchip.system.DefaultConfig.fir@224694.12]
  wire [3:0] _GEN_6909; // @[TLSimpleL2.scala 527:69:freechips.rocketchip.system.DefaultConfig.fir@224690.10]
  wire [3:0] _GEN_6910; // @[TLSimpleL2.scala 525:27:freechips.rocketchip.system.DefaultConfig.fir@224685.8]
  wire [3:0] _GEN_6912; // @[TLSimpleL2.scala 523:51:freechips.rocketchip.system.DefaultConfig.fir@224683.6]
  wire [3:0] _GEN_6922; // @[TLSimpleL2.scala 519:36:freechips.rocketchip.system.DefaultConfig.fir@224673.4]
  wire  _T_14102; // @[TLSimpleL2.scala 544:19:freechips.rocketchip.system.DefaultConfig.fir@224708.4]
  wire [2:0] _T_14104; // @[TLSimpleL2.scala 545:44:freechips.rocketchip.system.DefaultConfig.fir@224711.6]
  wire [3:0] _T_14106; // @[TLSimpleL2.scala 547:52:freechips.rocketchip.system.DefaultConfig.fir@224714.6]
  wire [2:0] _T_14107; // @[TLSimpleL2.scala 547:52:freechips.rocketchip.system.DefaultConfig.fir@224715.6]
  wire [7:0] _GEN_6924; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire [7:0] _GEN_6925; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire [7:0] _GEN_6926; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire [7:0] _GEN_6927; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire [7:0] _GEN_6928; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire [7:0] _GEN_6929; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire [7:0] _GEN_6930; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire  _T_14114; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  wire  _T_14115; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224717.6]
  wire  _T_14116; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224718.6]
  wire  _T_14117; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224719.6]
  wire  _T_14118; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224720.6]
  wire  _T_14119; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224721.6]
  wire  _T_14120; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224722.6]
  wire  _T_14121; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224723.6]
  wire [7:0] _T_14123; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224725.6]
  wire [7:0] _T_14125; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224727.6]
  wire [7:0] _T_14127; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224729.6]
  wire [7:0] _T_14129; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224731.6]
  wire [7:0] _T_14131; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224733.6]
  wire [7:0] _T_14133; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224735.6]
  wire [7:0] _T_14135; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224737.6]
  wire [7:0] _T_14137; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224739.6]
  wire [15:0] _T_14138; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224740.6]
  wire [15:0] _T_14139; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224741.6]
  wire [31:0] _T_14140; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224742.6]
  wire [15:0] _T_14141; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224743.6]
  wire [15:0] _T_14142; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224744.6]
  wire [31:0] _T_14143; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224745.6]
  wire [63:0] _T_14144; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224746.6]
  wire [63:0] _T_14145; // @[TLSimpleL2.scala 542:13:freechips.rocketchip.system.DefaultConfig.fir@224747.6]
  wire [63:0] _GEN_6932; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6933; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6934; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6935; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6936; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6937; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6938; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _T_14146; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  wire [63:0] _GEN_6940; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _GEN_6941; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _GEN_6942; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _GEN_6943; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _GEN_6944; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _GEN_6945; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _GEN_6946; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _T_14147; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  wire [63:0] _T_14148; // @[TLSimpleL2.scala 542:37:freechips.rocketchip.system.DefaultConfig.fir@224750.6]
  wire [3:0] _GEN_6955; // @[TLSimpleL2.scala 550:32:freechips.rocketchip.system.DefaultConfig.fir@224752.6]
  wire [3:0] _GEN_6965; // @[TLSimpleL2.scala 544:41:freechips.rocketchip.system.DefaultConfig.fir@224709.4]
  wire  _T_14151; // @[Counter.scala 34:24:freechips.rocketchip.system.DefaultConfig.fir@224759.6]
  wire [2:0] _T_14153; // @[Counter.scala 35:22:freechips.rocketchip.system.DefaultConfig.fir@224761.6]
  wire  _T_14154; // @[Counter.scala 64:20:freechips.rocketchip.system.DefaultConfig.fir@224764.4]
  wire  _T_14162; // @[TLSimpleL2.scala 562:36:freechips.rocketchip.system.DefaultConfig.fir@224773.4]
  wire [3:0] _GEN_6975; // @[TLSimpleL2.scala 563:20:freechips.rocketchip.system.DefaultConfig.fir@224775.6]
  wire [3:0] _GEN_6976; // @[TLSimpleL2.scala 562:51:freechips.rocketchip.system.DefaultConfig.fir@224774.4]
  wire [26:0] _T_14163; // @[TLSimpleL2.scala 574:30:freechips.rocketchip.system.DefaultConfig.fir@224782.4]
  wire [32:0] _T_14164; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224783.4]
  wire  _T_14268; // @[TLSimpleL2.scala 647:29:freechips.rocketchip.system.DefaultConfig.fir@224932.4]
  wire  _T_14269; // @[TLSimpleL2.scala 647:58:freechips.rocketchip.system.DefaultConfig.fir@224933.4]
  wire  _T_14270; // @[TLSimpleL2.scala 647:48:freechips.rocketchip.system.DefaultConfig.fir@224934.4]
  wire  _T_14168; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@224787.4]
  wire  _T_14170; // @[TLSimpleL2.scala 586:19:freechips.rocketchip.system.DefaultConfig.fir@224789.4]
  wire [3:0] _GEN_6977; // @[TLSimpleL2.scala 586:43:freechips.rocketchip.system.DefaultConfig.fir@224790.4]
  wire  _T_14172; // @[TLSimpleL2.scala 590:54:freechips.rocketchip.system.DefaultConfig.fir@224794.4]
  reg [2:0] value_2; // @[Counter.scala 26:33:freechips.rocketchip.system.DefaultConfig.fir@224795.4]
  reg [31:0] _RAND_2137;
  wire  _T_14174; // @[Counter.scala 34:24:freechips.rocketchip.system.DefaultConfig.fir@224797.6]
  wire [2:0] _T_14176; // @[Counter.scala 35:22:freechips.rocketchip.system.DefaultConfig.fir@224799.6]
  wire  _T_14177; // @[Counter.scala 64:20:freechips.rocketchip.system.DefaultConfig.fir@224802.4]
  wire  _T_14179; // @[TLSimpleL2.scala 591:38:freechips.rocketchip.system.DefaultConfig.fir@224804.4]
  wire [3:0] _GEN_6979; // @[TLSimpleL2.scala 591:50:freechips.rocketchip.system.DefaultConfig.fir@224805.4]
  wire  _T_14182; // @[TLSimpleL2.scala 597:40:freechips.rocketchip.system.DefaultConfig.fir@224810.4]
  wire  _T_14188; // @[TLSimpleL2.scala 612:42:freechips.rocketchip.system.DefaultConfig.fir@224827.4]
  wire  _T_14190; // @[TLSimpleL2.scala 615:62:freechips.rocketchip.system.DefaultConfig.fir@224832.4]
  reg [2:0] value_3; // @[Counter.scala 26:33:freechips.rocketchip.system.DefaultConfig.fir@224833.4]
  reg [31:0] _RAND_2138;
  wire  _T_14192; // @[Counter.scala 34:24:freechips.rocketchip.system.DefaultConfig.fir@224835.6]
  wire [2:0] _T_14194; // @[Counter.scala 35:22:freechips.rocketchip.system.DefaultConfig.fir@224837.6]
  wire  _T_14195; // @[Counter.scala 64:20:freechips.rocketchip.system.DefaultConfig.fir@224840.4]
  wire  _T_14197; // @[TLSimpleL2.scala 616:37:freechips.rocketchip.system.DefaultConfig.fir@224842.4]
  wire [63:0] _GEN_7004; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  wire [63:0] _GEN_7005; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  wire [63:0] _GEN_7006; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  wire [63:0] _GEN_7007; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  wire [63:0] _GEN_7008; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  wire [63:0] _GEN_7009; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  wire  _T_14272; // @[TLSimpleL2.scala 652:35:freechips.rocketchip.system.DefaultConfig.fir@224937.4]
  wire [2:0] _T_14274; // @[TLSimpleL2.scala 653:42:freechips.rocketchip.system.DefaultConfig.fir@224940.6]
  wire [3:0] _T_14283; // @[TLSimpleL2.scala 661:64:freechips.rocketchip.system.DefaultConfig.fir@224949.4]
  wire [2:0] _T_14284; // @[TLSimpleL2.scala 661:64:freechips.rocketchip.system.DefaultConfig.fir@224950.4]
  wire [63:0] _GEN_7015; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  wire [63:0] _GEN_7016; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  wire [63:0] _GEN_7017; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  wire [63:0] _GEN_7018; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  wire [63:0] _GEN_7019; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  wire [63:0] _GEN_7020; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  wire  _GEN_7033; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  wire  _GEN_7034; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  wire  _GEN_7035; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  wire  _GEN_7036; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  wire  _GEN_7041; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  wire  _GEN_7042; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  wire  _GEN_7043; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  wire  _GEN_7044; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  wire  _GEN_7049; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224190.10]
  wire  _GEN_7051; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7052; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7053; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7054; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7055; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7056; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7057; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  wire  _GEN_7066; // @[TLSimpleL2.scala 602:17:freechips.rocketchip.system.DefaultConfig.fir@224821.10]
  TLMonitor_54 TLMonitor ( // @[Nodes.scala 25:25:freechips.rocketchip.system.DefaultConfig.fir@220967.4]
    .clock(TLMonitor_clock),
    .reset(TLMonitor_reset),
    .io_in_a_ready(TLMonitor_io_in_a_ready),
    .io_in_a_valid(TLMonitor_io_in_a_valid),
    .io_in_a_bits_opcode(TLMonitor_io_in_a_bits_opcode),
    .io_in_a_bits_param(TLMonitor_io_in_a_bits_param),
    .io_in_a_bits_size(TLMonitor_io_in_a_bits_size),
    .io_in_a_bits_source(TLMonitor_io_in_a_bits_source),
    .io_in_a_bits_address(TLMonitor_io_in_a_bits_address),
    .io_in_a_bits_mask(TLMonitor_io_in_a_bits_mask),
    .io_in_a_bits_corrupt(TLMonitor_io_in_a_bits_corrupt),
    .io_in_d_ready(TLMonitor_io_in_d_ready),
    .io_in_d_valid(TLMonitor_io_in_d_valid),
    .io_in_d_bits_opcode(TLMonitor_io_in_d_bits_opcode),
    .io_in_d_bits_size(TLMonitor_io_in_d_bits_size),
    .io_in_d_bits_source(TLMonitor_io_in_d_bits_source)
  );
  L2_meta_array L2_meta_array ( // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@221200.4]
    .RW0_addr(L2_meta_array_RW0_addr),
    .RW0_en(L2_meta_array_RW0_en),
    .RW0_clk(L2_meta_array_RW0_clk),
    .RW0_wmode(L2_meta_array_RW0_wmode),
    .RW0_wdata_0_valid(L2_meta_array_RW0_wdata_0_valid),
    .RW0_wdata_0_dirty(L2_meta_array_RW0_wdata_0_dirty),
    .RW0_wdata_0_tag(L2_meta_array_RW0_wdata_0_tag),
    .RW0_wdata_0_rr_state(L2_meta_array_RW0_wdata_0_rr_state),
    .RW0_wdata_0_dsid(L2_meta_array_RW0_wdata_0_dsid),
    .RW0_wdata_1_valid(L2_meta_array_RW0_wdata_1_valid),
    .RW0_wdata_1_dirty(L2_meta_array_RW0_wdata_1_dirty),
    .RW0_wdata_1_tag(L2_meta_array_RW0_wdata_1_tag),
    .RW0_wdata_1_rr_state(L2_meta_array_RW0_wdata_1_rr_state),
    .RW0_wdata_1_dsid(L2_meta_array_RW0_wdata_1_dsid),
    .RW0_wdata_2_valid(L2_meta_array_RW0_wdata_2_valid),
    .RW0_wdata_2_dirty(L2_meta_array_RW0_wdata_2_dirty),
    .RW0_wdata_2_tag(L2_meta_array_RW0_wdata_2_tag),
    .RW0_wdata_2_rr_state(L2_meta_array_RW0_wdata_2_rr_state),
    .RW0_wdata_2_dsid(L2_meta_array_RW0_wdata_2_dsid),
    .RW0_wdata_3_valid(L2_meta_array_RW0_wdata_3_valid),
    .RW0_wdata_3_dirty(L2_meta_array_RW0_wdata_3_dirty),
    .RW0_wdata_3_tag(L2_meta_array_RW0_wdata_3_tag),
    .RW0_wdata_3_rr_state(L2_meta_array_RW0_wdata_3_rr_state),
    .RW0_wdata_3_dsid(L2_meta_array_RW0_wdata_3_dsid),
    .RW0_wdata_4_valid(L2_meta_array_RW0_wdata_4_valid),
    .RW0_wdata_4_dirty(L2_meta_array_RW0_wdata_4_dirty),
    .RW0_wdata_4_tag(L2_meta_array_RW0_wdata_4_tag),
    .RW0_wdata_4_rr_state(L2_meta_array_RW0_wdata_4_rr_state),
    .RW0_wdata_4_dsid(L2_meta_array_RW0_wdata_4_dsid),
    .RW0_wdata_5_valid(L2_meta_array_RW0_wdata_5_valid),
    .RW0_wdata_5_dirty(L2_meta_array_RW0_wdata_5_dirty),
    .RW0_wdata_5_tag(L2_meta_array_RW0_wdata_5_tag),
    .RW0_wdata_5_rr_state(L2_meta_array_RW0_wdata_5_rr_state),
    .RW0_wdata_5_dsid(L2_meta_array_RW0_wdata_5_dsid),
    .RW0_wdata_6_valid(L2_meta_array_RW0_wdata_6_valid),
    .RW0_wdata_6_dirty(L2_meta_array_RW0_wdata_6_dirty),
    .RW0_wdata_6_tag(L2_meta_array_RW0_wdata_6_tag),
    .RW0_wdata_6_rr_state(L2_meta_array_RW0_wdata_6_rr_state),
    .RW0_wdata_6_dsid(L2_meta_array_RW0_wdata_6_dsid),
    .RW0_wdata_7_valid(L2_meta_array_RW0_wdata_7_valid),
    .RW0_wdata_7_dirty(L2_meta_array_RW0_wdata_7_dirty),
    .RW0_wdata_7_tag(L2_meta_array_RW0_wdata_7_tag),
    .RW0_wdata_7_rr_state(L2_meta_array_RW0_wdata_7_rr_state),
    .RW0_wdata_7_dsid(L2_meta_array_RW0_wdata_7_dsid),
    .RW0_wdata_8_valid(L2_meta_array_RW0_wdata_8_valid),
    .RW0_wdata_8_dirty(L2_meta_array_RW0_wdata_8_dirty),
    .RW0_wdata_8_tag(L2_meta_array_RW0_wdata_8_tag),
    .RW0_wdata_8_rr_state(L2_meta_array_RW0_wdata_8_rr_state),
    .RW0_wdata_8_dsid(L2_meta_array_RW0_wdata_8_dsid),
    .RW0_wdata_9_valid(L2_meta_array_RW0_wdata_9_valid),
    .RW0_wdata_9_dirty(L2_meta_array_RW0_wdata_9_dirty),
    .RW0_wdata_9_tag(L2_meta_array_RW0_wdata_9_tag),
    .RW0_wdata_9_rr_state(L2_meta_array_RW0_wdata_9_rr_state),
    .RW0_wdata_9_dsid(L2_meta_array_RW0_wdata_9_dsid),
    .RW0_wdata_10_valid(L2_meta_array_RW0_wdata_10_valid),
    .RW0_wdata_10_dirty(L2_meta_array_RW0_wdata_10_dirty),
    .RW0_wdata_10_tag(L2_meta_array_RW0_wdata_10_tag),
    .RW0_wdata_10_rr_state(L2_meta_array_RW0_wdata_10_rr_state),
    .RW0_wdata_10_dsid(L2_meta_array_RW0_wdata_10_dsid),
    .RW0_wdata_11_valid(L2_meta_array_RW0_wdata_11_valid),
    .RW0_wdata_11_dirty(L2_meta_array_RW0_wdata_11_dirty),
    .RW0_wdata_11_tag(L2_meta_array_RW0_wdata_11_tag),
    .RW0_wdata_11_rr_state(L2_meta_array_RW0_wdata_11_rr_state),
    .RW0_wdata_11_dsid(L2_meta_array_RW0_wdata_11_dsid),
    .RW0_wdata_12_valid(L2_meta_array_RW0_wdata_12_valid),
    .RW0_wdata_12_dirty(L2_meta_array_RW0_wdata_12_dirty),
    .RW0_wdata_12_tag(L2_meta_array_RW0_wdata_12_tag),
    .RW0_wdata_12_rr_state(L2_meta_array_RW0_wdata_12_rr_state),
    .RW0_wdata_12_dsid(L2_meta_array_RW0_wdata_12_dsid),
    .RW0_wdata_13_valid(L2_meta_array_RW0_wdata_13_valid),
    .RW0_wdata_13_dirty(L2_meta_array_RW0_wdata_13_dirty),
    .RW0_wdata_13_tag(L2_meta_array_RW0_wdata_13_tag),
    .RW0_wdata_13_rr_state(L2_meta_array_RW0_wdata_13_rr_state),
    .RW0_wdata_13_dsid(L2_meta_array_RW0_wdata_13_dsid),
    .RW0_wdata_14_valid(L2_meta_array_RW0_wdata_14_valid),
    .RW0_wdata_14_dirty(L2_meta_array_RW0_wdata_14_dirty),
    .RW0_wdata_14_tag(L2_meta_array_RW0_wdata_14_tag),
    .RW0_wdata_14_rr_state(L2_meta_array_RW0_wdata_14_rr_state),
    .RW0_wdata_14_dsid(L2_meta_array_RW0_wdata_14_dsid),
    .RW0_wdata_15_valid(L2_meta_array_RW0_wdata_15_valid),
    .RW0_wdata_15_dirty(L2_meta_array_RW0_wdata_15_dirty),
    .RW0_wdata_15_tag(L2_meta_array_RW0_wdata_15_tag),
    .RW0_wdata_15_rr_state(L2_meta_array_RW0_wdata_15_rr_state),
    .RW0_wdata_15_dsid(L2_meta_array_RW0_wdata_15_dsid),
    .RW0_rdata_0_valid(L2_meta_array_RW0_rdata_0_valid),
    .RW0_rdata_0_dirty(L2_meta_array_RW0_rdata_0_dirty),
    .RW0_rdata_0_tag(L2_meta_array_RW0_rdata_0_tag),
    .RW0_rdata_0_rr_state(L2_meta_array_RW0_rdata_0_rr_state),
    .RW0_rdata_0_dsid(L2_meta_array_RW0_rdata_0_dsid),
    .RW0_rdata_1_valid(L2_meta_array_RW0_rdata_1_valid),
    .RW0_rdata_1_dirty(L2_meta_array_RW0_rdata_1_dirty),
    .RW0_rdata_1_tag(L2_meta_array_RW0_rdata_1_tag),
    .RW0_rdata_1_rr_state(L2_meta_array_RW0_rdata_1_rr_state),
    .RW0_rdata_1_dsid(L2_meta_array_RW0_rdata_1_dsid),
    .RW0_rdata_2_valid(L2_meta_array_RW0_rdata_2_valid),
    .RW0_rdata_2_dirty(L2_meta_array_RW0_rdata_2_dirty),
    .RW0_rdata_2_tag(L2_meta_array_RW0_rdata_2_tag),
    .RW0_rdata_2_rr_state(L2_meta_array_RW0_rdata_2_rr_state),
    .RW0_rdata_2_dsid(L2_meta_array_RW0_rdata_2_dsid),
    .RW0_rdata_3_valid(L2_meta_array_RW0_rdata_3_valid),
    .RW0_rdata_3_dirty(L2_meta_array_RW0_rdata_3_dirty),
    .RW0_rdata_3_tag(L2_meta_array_RW0_rdata_3_tag),
    .RW0_rdata_3_rr_state(L2_meta_array_RW0_rdata_3_rr_state),
    .RW0_rdata_3_dsid(L2_meta_array_RW0_rdata_3_dsid),
    .RW0_rdata_4_valid(L2_meta_array_RW0_rdata_4_valid),
    .RW0_rdata_4_dirty(L2_meta_array_RW0_rdata_4_dirty),
    .RW0_rdata_4_tag(L2_meta_array_RW0_rdata_4_tag),
    .RW0_rdata_4_rr_state(L2_meta_array_RW0_rdata_4_rr_state),
    .RW0_rdata_4_dsid(L2_meta_array_RW0_rdata_4_dsid),
    .RW0_rdata_5_valid(L2_meta_array_RW0_rdata_5_valid),
    .RW0_rdata_5_dirty(L2_meta_array_RW0_rdata_5_dirty),
    .RW0_rdata_5_tag(L2_meta_array_RW0_rdata_5_tag),
    .RW0_rdata_5_rr_state(L2_meta_array_RW0_rdata_5_rr_state),
    .RW0_rdata_5_dsid(L2_meta_array_RW0_rdata_5_dsid),
    .RW0_rdata_6_valid(L2_meta_array_RW0_rdata_6_valid),
    .RW0_rdata_6_dirty(L2_meta_array_RW0_rdata_6_dirty),
    .RW0_rdata_6_tag(L2_meta_array_RW0_rdata_6_tag),
    .RW0_rdata_6_rr_state(L2_meta_array_RW0_rdata_6_rr_state),
    .RW0_rdata_6_dsid(L2_meta_array_RW0_rdata_6_dsid),
    .RW0_rdata_7_valid(L2_meta_array_RW0_rdata_7_valid),
    .RW0_rdata_7_dirty(L2_meta_array_RW0_rdata_7_dirty),
    .RW0_rdata_7_tag(L2_meta_array_RW0_rdata_7_tag),
    .RW0_rdata_7_rr_state(L2_meta_array_RW0_rdata_7_rr_state),
    .RW0_rdata_7_dsid(L2_meta_array_RW0_rdata_7_dsid),
    .RW0_rdata_8_valid(L2_meta_array_RW0_rdata_8_valid),
    .RW0_rdata_8_dirty(L2_meta_array_RW0_rdata_8_dirty),
    .RW0_rdata_8_tag(L2_meta_array_RW0_rdata_8_tag),
    .RW0_rdata_8_rr_state(L2_meta_array_RW0_rdata_8_rr_state),
    .RW0_rdata_8_dsid(L2_meta_array_RW0_rdata_8_dsid),
    .RW0_rdata_9_valid(L2_meta_array_RW0_rdata_9_valid),
    .RW0_rdata_9_dirty(L2_meta_array_RW0_rdata_9_dirty),
    .RW0_rdata_9_tag(L2_meta_array_RW0_rdata_9_tag),
    .RW0_rdata_9_rr_state(L2_meta_array_RW0_rdata_9_rr_state),
    .RW0_rdata_9_dsid(L2_meta_array_RW0_rdata_9_dsid),
    .RW0_rdata_10_valid(L2_meta_array_RW0_rdata_10_valid),
    .RW0_rdata_10_dirty(L2_meta_array_RW0_rdata_10_dirty),
    .RW0_rdata_10_tag(L2_meta_array_RW0_rdata_10_tag),
    .RW0_rdata_10_rr_state(L2_meta_array_RW0_rdata_10_rr_state),
    .RW0_rdata_10_dsid(L2_meta_array_RW0_rdata_10_dsid),
    .RW0_rdata_11_valid(L2_meta_array_RW0_rdata_11_valid),
    .RW0_rdata_11_dirty(L2_meta_array_RW0_rdata_11_dirty),
    .RW0_rdata_11_tag(L2_meta_array_RW0_rdata_11_tag),
    .RW0_rdata_11_rr_state(L2_meta_array_RW0_rdata_11_rr_state),
    .RW0_rdata_11_dsid(L2_meta_array_RW0_rdata_11_dsid),
    .RW0_rdata_12_valid(L2_meta_array_RW0_rdata_12_valid),
    .RW0_rdata_12_dirty(L2_meta_array_RW0_rdata_12_dirty),
    .RW0_rdata_12_tag(L2_meta_array_RW0_rdata_12_tag),
    .RW0_rdata_12_rr_state(L2_meta_array_RW0_rdata_12_rr_state),
    .RW0_rdata_12_dsid(L2_meta_array_RW0_rdata_12_dsid),
    .RW0_rdata_13_valid(L2_meta_array_RW0_rdata_13_valid),
    .RW0_rdata_13_dirty(L2_meta_array_RW0_rdata_13_dirty),
    .RW0_rdata_13_tag(L2_meta_array_RW0_rdata_13_tag),
    .RW0_rdata_13_rr_state(L2_meta_array_RW0_rdata_13_rr_state),
    .RW0_rdata_13_dsid(L2_meta_array_RW0_rdata_13_dsid),
    .RW0_rdata_14_valid(L2_meta_array_RW0_rdata_14_valid),
    .RW0_rdata_14_dirty(L2_meta_array_RW0_rdata_14_dirty),
    .RW0_rdata_14_tag(L2_meta_array_RW0_rdata_14_tag),
    .RW0_rdata_14_rr_state(L2_meta_array_RW0_rdata_14_rr_state),
    .RW0_rdata_14_dsid(L2_meta_array_RW0_rdata_14_dsid),
    .RW0_rdata_15_valid(L2_meta_array_RW0_rdata_15_valid),
    .RW0_rdata_15_dirty(L2_meta_array_RW0_rdata_15_dirty),
    .RW0_rdata_15_tag(L2_meta_array_RW0_rdata_15_tag),
    .RW0_rdata_15_rr_state(L2_meta_array_RW0_rdata_15_rr_state),
    .RW0_rdata_15_dsid(L2_meta_array_RW0_rdata_15_dsid)
  );
  L2_data_array L2_data_array ( // @[DescribedSRAM.scala 23:21:freechips.rocketchip.system.DefaultConfig.fir@224556.4]
    .RW0_addr(L2_data_array_RW0_addr),
    .RW0_en(L2_data_array_RW0_en),
    .RW0_clk(L2_data_array_RW0_clk),
    .RW0_wmode(L2_data_array_RW0_wmode),
    .RW0_wdata_0(L2_data_array_RW0_wdata_0),
    .RW0_wdata_1(L2_data_array_RW0_wdata_1),
    .RW0_wdata_2(L2_data_array_RW0_wdata_2),
    .RW0_wdata_3(L2_data_array_RW0_wdata_3),
    .RW0_wdata_4(L2_data_array_RW0_wdata_4),
    .RW0_wdata_5(L2_data_array_RW0_wdata_5),
    .RW0_wdata_6(L2_data_array_RW0_wdata_6),
    .RW0_wdata_7(L2_data_array_RW0_wdata_7),
    .RW0_wdata_8(L2_data_array_RW0_wdata_8),
    .RW0_wdata_9(L2_data_array_RW0_wdata_9),
    .RW0_wdata_10(L2_data_array_RW0_wdata_10),
    .RW0_wdata_11(L2_data_array_RW0_wdata_11),
    .RW0_wdata_12(L2_data_array_RW0_wdata_12),
    .RW0_wdata_13(L2_data_array_RW0_wdata_13),
    .RW0_wdata_14(L2_data_array_RW0_wdata_14),
    .RW0_wdata_15(L2_data_array_RW0_wdata_15),
    .RW0_rdata_0(L2_data_array_RW0_rdata_0),
    .RW0_rdata_1(L2_data_array_RW0_rdata_1),
    .RW0_rdata_2(L2_data_array_RW0_rdata_2),
    .RW0_rdata_3(L2_data_array_RW0_rdata_3),
    .RW0_rdata_4(L2_data_array_RW0_rdata_4),
    .RW0_rdata_5(L2_data_array_RW0_rdata_5),
    .RW0_rdata_6(L2_data_array_RW0_rdata_6),
    .RW0_rdata_7(L2_data_array_RW0_rdata_7),
    .RW0_rdata_8(L2_data_array_RW0_rdata_8),
    .RW0_rdata_9(L2_data_array_RW0_rdata_9),
    .RW0_rdata_10(L2_data_array_RW0_rdata_10),
    .RW0_rdata_11(L2_data_array_RW0_rdata_11),
    .RW0_rdata_12(L2_data_array_RW0_rdata_12),
    .RW0_rdata_13(L2_data_array_RW0_rdata_13),
    .RW0_rdata_14(L2_data_array_RW0_rdata_14),
    .RW0_rdata_15(L2_data_array_RW0_rdata_15),
    .RW0_wmask_0(L2_data_array_RW0_wmask_0),
    .RW0_wmask_1(L2_data_array_RW0_wmask_1),
    .RW0_wmask_2(L2_data_array_RW0_wmask_2),
    .RW0_wmask_3(L2_data_array_RW0_wmask_3),
    .RW0_wmask_4(L2_data_array_RW0_wmask_4),
    .RW0_wmask_5(L2_data_array_RW0_wmask_5),
    .RW0_wmask_6(L2_data_array_RW0_wmask_6),
    .RW0_wmask_7(L2_data_array_RW0_wmask_7),
    .RW0_wmask_8(L2_data_array_RW0_wmask_8),
    .RW0_wmask_9(L2_data_array_RW0_wmask_9),
    .RW0_wmask_10(L2_data_array_RW0_wmask_10),
    .RW0_wmask_11(L2_data_array_RW0_wmask_11),
    .RW0_wmask_12(L2_data_array_RW0_wmask_12),
    .RW0_wmask_13(L2_data_array_RW0_wmask_13),
    .RW0_wmask_14(L2_data_array_RW0_wmask_14),
    .RW0_wmask_15(L2_data_array_RW0_wmask_15)
  );
  assign _T_259 = _T_258 < 13'h1000; // @[TLSimpleL2.scala 90:26:freechips.rocketchip.system.DefaultConfig.fir@221009.4]
  assign _T_261 = reset == 1'h0; // @[TLSimpleL2.scala 90:48:freechips.rocketchip.system.DefaultConfig.fir@221011.4]
  assign _T_262 = _T_259 & _T_261; // @[TLSimpleL2.scala 90:45:freechips.rocketchip.system.DefaultConfig.fir@221012.4]
  assign _T_264 = _T_258 + 13'h1; // @[TLSimpleL2.scala 91:39:freechips.rocketchip.system.DefaultConfig.fir@221015.6]
  assign _T_335 = _T_267 == 4'h0; // @[TLSimpleL2.scala 243:36:freechips.rocketchip.system.DefaultConfig.fir@221121.4]
  assign _T_336 = _T_262 == 1'h0; // @[TLSimpleL2.scala 243:50:freechips.rocketchip.system.DefaultConfig.fir@221122.4]
  assign _T_337 = _T_335 & _T_336; // @[TLSimpleL2.scala 243:47:freechips.rocketchip.system.DefaultConfig.fir@221123.4]
  assign _T_451 = _T_337 | _T_337; // @[TLSimpleL2.scala 272:45:freechips.rocketchip.system.DefaultConfig.fir@221188.4]
  assign _T_426 = _T_267 == 4'h1; // @[TLSimpleL2.scala 250:36:freechips.rocketchip.system.DefaultConfig.fir@221147.4]
  assign _T_452 = _T_451 | _T_426; // @[TLSimpleL2.scala 272:65:freechips.rocketchip.system.DefaultConfig.fir@221189.4]
  assign _T_273 = _T_452 & auto_in_a_valid; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@221030.4]
  assign _T_14180 = _T_267 == 4'hb; // @[TLSimpleL2.scala 595:35:freechips.rocketchip.system.DefaultConfig.fir@224808.4]
  assign _T_14199 = _T_267 == 4'hd; // @[TLSimpleL2.scala 627:34:freechips.rocketchip.system.DefaultConfig.fir@224854.4]
  assign _T_14267 = _T_14180 | _T_14199; // @[TLSimpleL2.scala 644:38:freechips.rocketchip.system.DefaultConfig.fir@224930.4]
  assign _T_274 = auto_out_a_ready & _T_14267; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@221033.4]
  assign _T_275 = auto_in_a_bits_size >= 3'h3; // @[TLSimpleL2.scala 168:41:freechips.rocketchip.system.DefaultConfig.fir@221036.4]
  assign _T_276 = 8'h1 << auto_in_a_bits_size; // @[TLSimpleL2.scala 169:45:freechips.rocketchip.system.DefaultConfig.fir@221037.4]
  assign _T_277 = _T_276[7:3]; // @[TLSimpleL2.scala 169:64:freechips.rocketchip.system.DefaultConfig.fir@221038.4]
  assign _T_278 = _T_277 - 5'h1; // @[TLSimpleL2.scala 169:82:freechips.rocketchip.system.DefaultConfig.fir@221039.4]
  assign _T_279 = $unsigned(_T_278); // @[TLSimpleL2.scala 169:82:freechips.rocketchip.system.DefaultConfig.fir@221040.4]
  assign _T_280 = _T_279[4:0]; // @[TLSimpleL2.scala 169:82:freechips.rocketchip.system.DefaultConfig.fir@221041.4]
  assign _T_281 = _T_275 ? _T_280 : 5'h0; // @[TLSimpleL2.scala 169:24:freechips.rocketchip.system.DefaultConfig.fir@221042.4]
  assign _T_283 = auto_in_a_bits_opcode == 3'h4; // @[TLSimpleL2.scala 174:52:freechips.rocketchip.system.DefaultConfig.fir@221044.4]
  assign _T_284 = _T_273 & _T_283; // @[TLSimpleL2.scala 174:38:freechips.rocketchip.system.DefaultConfig.fir@221045.4]
  assign _T_285 = auto_in_a_bits_opcode == 3'h0; // @[TLSimpleL2.scala 175:53:freechips.rocketchip.system.DefaultConfig.fir@221046.4]
  assign _T_286 = auto_in_a_bits_opcode == 3'h1; // @[TLSimpleL2.scala 175:93:freechips.rocketchip.system.DefaultConfig.fir@221047.4]
  assign _T_287 = _T_285 | _T_286; // @[TLSimpleL2.scala 175:80:freechips.rocketchip.system.DefaultConfig.fir@221048.4]
  assign _T_288 = _T_273 & _T_287; // @[TLSimpleL2.scala 175:39:freechips.rocketchip.system.DefaultConfig.fir@221049.4]
  assign _T_456 = _T_267 == 4'h2; // @[TLSimpleL2.scala 279:31:freechips.rocketchip.system.DefaultConfig.fir@221194.4]
  assign _T_14286 = _T_267 == 4'hf; // @[TLSimpleL2.scala 664:30:freechips.rocketchip.system.DefaultConfig.fir@224952.4]
  assign _T_14287 = _T_456 | _T_14286; // @[TLSimpleL2.scala 666:33:freechips.rocketchip.system.DefaultConfig.fir@224953.4]
  assign _T_289 = auto_in_d_ready & _T_14287; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@221050.4]
  assign _T_304 = auto_in_a_bits_address[5:3]; // @[TLSimpleL2.scala 191:31:freechips.rocketchip.system.DefaultConfig.fir@221058.4]
  assign _GEN_7022 = {{2'd0}, _T_304}; // @[TLSimpleL2.scala 193:61:freechips.rocketchip.system.DefaultConfig.fir@221061.4]
  assign _T_309 = _GEN_7022 + _T_281; // @[TLSimpleL2.scala 193:61:freechips.rocketchip.system.DefaultConfig.fir@221062.4]
  assign _T_310 = _T_335 ? _T_309 : {{1'd0}, _T_306}; // @[TLSimpleL2.scala 193:31:freechips.rocketchip.system.DefaultConfig.fir@221063.4]
  assign _T_314 = _T_335 ? _T_304 : _T_312; // @[TLSimpleL2.scala 195:33:freechips.rocketchip.system.DefaultConfig.fir@221066.4]
  assign _GEN_7023 = {{2'd0}, _T_314}; // @[TLSimpleL2.scala 196:47:freechips.rocketchip.system.DefaultConfig.fir@221067.4]
  assign _T_315 = _GEN_7023 == _T_310; // @[TLSimpleL2.scala 196:47:freechips.rocketchip.system.DefaultConfig.fir@221067.4]
  assign _GEN_7024 = {{2'd0}, _T_317}; // @[TLSimpleL2.scala 198:45:freechips.rocketchip.system.DefaultConfig.fir@221069.4]
  assign _T_318 = _GEN_7024 == _T_310; // @[TLSimpleL2.scala 198:45:freechips.rocketchip.system.DefaultConfig.fir@221069.4]
  assign _GEN_7025 = {{2'd0}, _T_320}; // @[TLSimpleL2.scala 200:43:freechips.rocketchip.system.DefaultConfig.fir@221071.4]
  assign _T_321 = _GEN_7025 == _T_310; // @[TLSimpleL2.scala 200:43:freechips.rocketchip.system.DefaultConfig.fir@221071.4]
  assign _GEN_8 = _T_288 ? auto_in_a_bits_dsid : {{1'd0}, _T_297}; // @[TLSimpleL2.scala 223:36:freechips.rocketchip.system.DefaultConfig.fir@221090.8]
  assign _GEN_12 = _T_288 ? _T_309 : {{1'd0}, _T_306}; // @[TLSimpleL2.scala 223:36:freechips.rocketchip.system.DefaultConfig.fir@221090.8]
  assign _GEN_13 = _T_288 ? 4'h1 : _T_267; // @[TLSimpleL2.scala 223:36:freechips.rocketchip.system.DefaultConfig.fir@221090.8]
  assign _GEN_19 = _T_284 ? auto_in_a_bits_dsid : _GEN_8; // @[TLSimpleL2.scala 207:28:freechips.rocketchip.system.DefaultConfig.fir@221074.6]
  assign _GEN_23 = _T_284 ? _T_309 : _GEN_12; // @[TLSimpleL2.scala 207:28:freechips.rocketchip.system.DefaultConfig.fir@221074.6]
  assign _GEN_24 = _T_284 ? 4'h4 : _GEN_13; // @[TLSimpleL2.scala 207:28:freechips.rocketchip.system.DefaultConfig.fir@221074.6]
  assign _GEN_30 = _T_335 ? _GEN_19 : {{1'd0}, _T_297}; // @[TLSimpleL2.scala 206:31:freechips.rocketchip.system.DefaultConfig.fir@221073.4]
  assign _GEN_34 = _T_335 ? _GEN_23 : {{1'd0}, _T_306}; // @[TLSimpleL2.scala 206:31:freechips.rocketchip.system.DefaultConfig.fir@221073.4]
  assign _GEN_35 = _T_335 ? _GEN_24 : _T_267; // @[TLSimpleL2.scala 206:31:freechips.rocketchip.system.DefaultConfig.fir@221073.4]
  assign _T_428 = _T_426 & _T_273; // @[TLSimpleL2.scala 254:60:freechips.rocketchip.system.DefaultConfig.fir@221149.4]
  assign _T_429 = _T_288 | _T_428; // @[TLSimpleL2.scala 254:26:freechips.rocketchip.system.DefaultConfig.fir@221150.4]
  assign _T_432 = _T_304 + 3'h1; // @[TLSimpleL2.scala 256:46:freechips.rocketchip.system.DefaultConfig.fir@221155.8]
  assign _T_435 = _T_312 + 3'h1; // @[TLSimpleL2.scala 258:56:freechips.rocketchip.system.DefaultConfig.fir@221162.10]
  assign _T_440 = {{1'd0}, _T_314}; // @[TLSimpleL2.scala 264:56:freechips.rocketchip.system.DefaultConfig.fir@221175.6]
  assign _T_441 = _T_440[2:0]; // @[TLSimpleL2.scala 264:56:freechips.rocketchip.system.DefaultConfig.fir@221176.6]
  assign _GEN_54 = _T_315 ? 4'h2 : _GEN_35; // @[TLSimpleL2.scala 267:33:freechips.rocketchip.system.DefaultConfig.fir@221184.6]
  assign _GEN_72 = _T_429 ? _GEN_54 : _GEN_35; // @[TLSimpleL2.scala 254:78:freechips.rocketchip.system.DefaultConfig.fir@221151.4]
  assign _T_458 = _T_456 & _T_289; // @[TLSimpleL2.scala 281:36:freechips.rocketchip.system.DefaultConfig.fir@221196.4]
  assign _GEN_73 = _T_458 ? 4'h4 : _GEN_72; // @[TLSimpleL2.scala 281:51:freechips.rocketchip.system.DefaultConfig.fir@221197.4]
  assign _T_481 = _T_291[16:6]; // @[TLSimpleL2.scala 298:21:freechips.rocketchip.system.DefaultConfig.fir@221201.4]
  assign _T_482 = _T_267 == 4'h6; // @[TLSimpleL2.scala 300:41:freechips.rocketchip.system.DefaultConfig.fir@221202.4]
  assign _T_483 = _T_262 | _T_482; // @[TLSimpleL2.scala 300:32:freechips.rocketchip.system.DefaultConfig.fir@221203.4]
  assign _T_484 = _T_267 == 4'h4; // @[TLSimpleL2.scala 301:33:freechips.rocketchip.system.DefaultConfig.fir@221204.4]
  assign _T_485 = _T_483 == 1'h0; // @[TLSimpleL2.scala 302:61:freechips.rocketchip.system.DefaultConfig.fir@221205.4]
  assign _T_486 = _T_484 & _T_485; // @[TLSimpleL2.scala 302:58:freechips.rocketchip.system.DefaultConfig.fir@221206.4]
  assign _T_530_1 = L2_meta_array_RW0_rdata_1_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221219.4]
  assign _T_530_0 = L2_meta_array_RW0_rdata_0_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221218.4]
  assign _T_549 = {_T_530_1,_T_530_0}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221234.4]
  assign _T_530_3 = L2_meta_array_RW0_rdata_3_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221221.4]
  assign _T_530_2 = L2_meta_array_RW0_rdata_2_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221220.4]
  assign _T_550 = {_T_530_3,_T_530_2}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221235.4]
  assign _T_551 = {_T_550,_T_549}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221236.4]
  assign _T_530_5 = L2_meta_array_RW0_rdata_5_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221223.4]
  assign _T_530_4 = L2_meta_array_RW0_rdata_4_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221222.4]
  assign _T_552 = {_T_530_5,_T_530_4}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221237.4]
  assign _T_530_7 = L2_meta_array_RW0_rdata_7_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221225.4]
  assign _T_530_6 = L2_meta_array_RW0_rdata_6_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221224.4]
  assign _T_553 = {_T_530_7,_T_530_6}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221238.4]
  assign _T_554 = {_T_553,_T_552}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221239.4]
  assign _T_555 = {_T_554,_T_551}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221240.4]
  assign _T_530_9 = L2_meta_array_RW0_rdata_9_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221227.4]
  assign _T_530_8 = L2_meta_array_RW0_rdata_8_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221226.4]
  assign _T_556 = {_T_530_9,_T_530_8}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221241.4]
  assign _T_530_11 = L2_meta_array_RW0_rdata_11_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221229.4]
  assign _T_530_10 = L2_meta_array_RW0_rdata_10_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221228.4]
  assign _T_557 = {_T_530_11,_T_530_10}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221242.4]
  assign _T_558 = {_T_557,_T_556}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221243.4]
  assign _T_530_13 = L2_meta_array_RW0_rdata_13_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221231.4]
  assign _T_530_12 = L2_meta_array_RW0_rdata_12_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221230.4]
  assign _T_559 = {_T_530_13,_T_530_12}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221244.4]
  assign _T_530_15 = L2_meta_array_RW0_rdata_15_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221233.4]
  assign _T_530_14 = L2_meta_array_RW0_rdata_14_valid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221216.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221232.4]
  assign _T_560 = {_T_530_15,_T_530_14}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221245.4]
  assign _T_561 = {_T_560,_T_559}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221246.4]
  assign _T_562 = {_T_561,_T_558}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221247.4]
  assign _T_563 = {_T_562,_T_555}; // @[TLSimpleL2.scala 306:62:freechips.rocketchip.system.DefaultConfig.fir@221248.4]
  assign _T_567_1 = L2_meta_array_RW0_rdata_1_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221252.4]
  assign _T_567_0 = L2_meta_array_RW0_rdata_0_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221251.4]
  assign _T_586 = {_T_567_1,_T_567_0}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221267.4]
  assign _T_567_3 = L2_meta_array_RW0_rdata_3_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221254.4]
  assign _T_567_2 = L2_meta_array_RW0_rdata_2_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221253.4]
  assign _T_587 = {_T_567_3,_T_567_2}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221268.4]
  assign _T_588 = {_T_587,_T_586}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221269.4]
  assign _T_567_5 = L2_meta_array_RW0_rdata_5_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221256.4]
  assign _T_567_4 = L2_meta_array_RW0_rdata_4_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221255.4]
  assign _T_589 = {_T_567_5,_T_567_4}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221270.4]
  assign _T_567_7 = L2_meta_array_RW0_rdata_7_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221258.4]
  assign _T_567_6 = L2_meta_array_RW0_rdata_6_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221257.4]
  assign _T_590 = {_T_567_7,_T_567_6}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221271.4]
  assign _T_591 = {_T_590,_T_589}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221272.4]
  assign _T_592 = {_T_591,_T_588}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221273.4]
  assign _T_567_9 = L2_meta_array_RW0_rdata_9_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221260.4]
  assign _T_567_8 = L2_meta_array_RW0_rdata_8_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221259.4]
  assign _T_593 = {_T_567_9,_T_567_8}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221274.4]
  assign _T_567_11 = L2_meta_array_RW0_rdata_11_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221262.4]
  assign _T_567_10 = L2_meta_array_RW0_rdata_10_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221261.4]
  assign _T_594 = {_T_567_11,_T_567_10}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221275.4]
  assign _T_595 = {_T_594,_T_593}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221276.4]
  assign _T_567_13 = L2_meta_array_RW0_rdata_13_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221264.4]
  assign _T_567_12 = L2_meta_array_RW0_rdata_12_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221263.4]
  assign _T_596 = {_T_567_13,_T_567_12}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221277.4]
  assign _T_567_15 = L2_meta_array_RW0_rdata_15_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221266.4]
  assign _T_567_14 = L2_meta_array_RW0_rdata_14_dirty; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221249.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221265.4]
  assign _T_597 = {_T_567_15,_T_567_14}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221278.4]
  assign _T_598 = {_T_597,_T_596}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221279.4]
  assign _T_599 = {_T_598,_T_595}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221280.4]
  assign _T_600 = {_T_599,_T_592}; // @[TLSimpleL2.scala 307:62:freechips.rocketchip.system.DefaultConfig.fir@221281.4]
  assign _T_626_1 = L2_meta_array_RW0_rdata_1_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221303.4]
  assign _T_626_0 = L2_meta_array_RW0_rdata_0_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221302.4]
  assign _T_645 = {_T_626_1,_T_626_0}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221318.4]
  assign _T_626_3 = L2_meta_array_RW0_rdata_3_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221305.4]
  assign _T_626_2 = L2_meta_array_RW0_rdata_2_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221304.4]
  assign _T_646 = {_T_626_3,_T_626_2}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221319.4]
  assign _T_647 = {_T_646,_T_645}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221320.4]
  assign _T_626_5 = L2_meta_array_RW0_rdata_5_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221307.4]
  assign _T_626_4 = L2_meta_array_RW0_rdata_4_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221306.4]
  assign _T_648 = {_T_626_5,_T_626_4}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221321.4]
  assign _T_626_7 = L2_meta_array_RW0_rdata_7_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221309.4]
  assign _T_626_6 = L2_meta_array_RW0_rdata_6_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221308.4]
  assign _T_649 = {_T_626_7,_T_626_6}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221322.4]
  assign _T_650 = {_T_649,_T_648}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221323.4]
  assign _T_651 = {_T_650,_T_647}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221324.4]
  assign _T_626_9 = L2_meta_array_RW0_rdata_9_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221311.4]
  assign _T_626_8 = L2_meta_array_RW0_rdata_8_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221310.4]
  assign _T_652 = {_T_626_9,_T_626_8}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221325.4]
  assign _T_626_11 = L2_meta_array_RW0_rdata_11_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221313.4]
  assign _T_626_10 = L2_meta_array_RW0_rdata_10_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221312.4]
  assign _T_653 = {_T_626_11,_T_626_10}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221326.4]
  assign _T_654 = {_T_653,_T_652}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221327.4]
  assign _T_626_13 = L2_meta_array_RW0_rdata_13_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221315.4]
  assign _T_626_12 = L2_meta_array_RW0_rdata_12_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221314.4]
  assign _T_655 = {_T_626_13,_T_626_12}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221328.4]
  assign _T_626_15 = L2_meta_array_RW0_rdata_15_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221317.4]
  assign _T_626_14 = L2_meta_array_RW0_rdata_14_rr_state; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221300.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221316.4]
  assign _T_656 = {_T_626_15,_T_626_14}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221329.4]
  assign _T_657 = {_T_656,_T_655}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221330.4]
  assign _T_658 = {_T_657,_T_654}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221331.4]
  assign _T_659 = {_T_658,_T_651}; // @[TLSimpleL2.scala 309:67:freechips.rocketchip.system.DefaultConfig.fir@221332.4]
  assign _GEN_78 = _T_484 ? 4'h5 : _GEN_73; // @[TLSimpleL2.scala 312:39:freechips.rocketchip.system.DefaultConfig.fir@221352.4]
  assign _T_13036 = _T_267 == 4'h5; // @[TLSimpleL2.scala 326:19:freechips.rocketchip.system.DefaultConfig.fir@223411.4]
  assign _GEN_80 = 11'h1 == _T_481 ? _T_6887_1 : _T_6887_0; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_81 = 11'h2 == _T_481 ? _T_6887_2 : _GEN_80; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_82 = 11'h3 == _T_481 ? _T_6887_3 : _GEN_81; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_83 = 11'h4 == _T_481 ? _T_6887_4 : _GEN_82; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_84 = 11'h5 == _T_481 ? _T_6887_5 : _GEN_83; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_85 = 11'h6 == _T_481 ? _T_6887_6 : _GEN_84; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_86 = 11'h7 == _T_481 ? _T_6887_7 : _GEN_85; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_87 = 11'h8 == _T_481 ? _T_6887_8 : _GEN_86; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_88 = 11'h9 == _T_481 ? _T_6887_9 : _GEN_87; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_89 = 11'ha == _T_481 ? _T_6887_10 : _GEN_88; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_90 = 11'hb == _T_481 ? _T_6887_11 : _GEN_89; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_91 = 11'hc == _T_481 ? _T_6887_12 : _GEN_90; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_92 = 11'hd == _T_481 ? _T_6887_13 : _GEN_91; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_93 = 11'he == _T_481 ? _T_6887_14 : _GEN_92; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_94 = 11'hf == _T_481 ? _T_6887_15 : _GEN_93; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_95 = 11'h10 == _T_481 ? _T_6887_16 : _GEN_94; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_96 = 11'h11 == _T_481 ? _T_6887_17 : _GEN_95; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_97 = 11'h12 == _T_481 ? _T_6887_18 : _GEN_96; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_98 = 11'h13 == _T_481 ? _T_6887_19 : _GEN_97; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_99 = 11'h14 == _T_481 ? _T_6887_20 : _GEN_98; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_100 = 11'h15 == _T_481 ? _T_6887_21 : _GEN_99; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_101 = 11'h16 == _T_481 ? _T_6887_22 : _GEN_100; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_102 = 11'h17 == _T_481 ? _T_6887_23 : _GEN_101; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_103 = 11'h18 == _T_481 ? _T_6887_24 : _GEN_102; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_104 = 11'h19 == _T_481 ? _T_6887_25 : _GEN_103; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_105 = 11'h1a == _T_481 ? _T_6887_26 : _GEN_104; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_106 = 11'h1b == _T_481 ? _T_6887_27 : _GEN_105; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_107 = 11'h1c == _T_481 ? _T_6887_28 : _GEN_106; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_108 = 11'h1d == _T_481 ? _T_6887_29 : _GEN_107; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_109 = 11'h1e == _T_481 ? _T_6887_30 : _GEN_108; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_110 = 11'h1f == _T_481 ? _T_6887_31 : _GEN_109; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_111 = 11'h20 == _T_481 ? _T_6887_32 : _GEN_110; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_112 = 11'h21 == _T_481 ? _T_6887_33 : _GEN_111; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_113 = 11'h22 == _T_481 ? _T_6887_34 : _GEN_112; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_114 = 11'h23 == _T_481 ? _T_6887_35 : _GEN_113; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_115 = 11'h24 == _T_481 ? _T_6887_36 : _GEN_114; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_116 = 11'h25 == _T_481 ? _T_6887_37 : _GEN_115; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_117 = 11'h26 == _T_481 ? _T_6887_38 : _GEN_116; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_118 = 11'h27 == _T_481 ? _T_6887_39 : _GEN_117; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_119 = 11'h28 == _T_481 ? _T_6887_40 : _GEN_118; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_120 = 11'h29 == _T_481 ? _T_6887_41 : _GEN_119; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_121 = 11'h2a == _T_481 ? _T_6887_42 : _GEN_120; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_122 = 11'h2b == _T_481 ? _T_6887_43 : _GEN_121; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_123 = 11'h2c == _T_481 ? _T_6887_44 : _GEN_122; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_124 = 11'h2d == _T_481 ? _T_6887_45 : _GEN_123; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_125 = 11'h2e == _T_481 ? _T_6887_46 : _GEN_124; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_126 = 11'h2f == _T_481 ? _T_6887_47 : _GEN_125; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_127 = 11'h30 == _T_481 ? _T_6887_48 : _GEN_126; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_128 = 11'h31 == _T_481 ? _T_6887_49 : _GEN_127; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_129 = 11'h32 == _T_481 ? _T_6887_50 : _GEN_128; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_130 = 11'h33 == _T_481 ? _T_6887_51 : _GEN_129; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_131 = 11'h34 == _T_481 ? _T_6887_52 : _GEN_130; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_132 = 11'h35 == _T_481 ? _T_6887_53 : _GEN_131; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_133 = 11'h36 == _T_481 ? _T_6887_54 : _GEN_132; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_134 = 11'h37 == _T_481 ? _T_6887_55 : _GEN_133; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_135 = 11'h38 == _T_481 ? _T_6887_56 : _GEN_134; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_136 = 11'h39 == _T_481 ? _T_6887_57 : _GEN_135; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_137 = 11'h3a == _T_481 ? _T_6887_58 : _GEN_136; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_138 = 11'h3b == _T_481 ? _T_6887_59 : _GEN_137; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_139 = 11'h3c == _T_481 ? _T_6887_60 : _GEN_138; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_140 = 11'h3d == _T_481 ? _T_6887_61 : _GEN_139; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_141 = 11'h3e == _T_481 ? _T_6887_62 : _GEN_140; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_142 = 11'h3f == _T_481 ? _T_6887_63 : _GEN_141; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_143 = 11'h40 == _T_481 ? _T_6887_64 : _GEN_142; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_144 = 11'h41 == _T_481 ? _T_6887_65 : _GEN_143; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_145 = 11'h42 == _T_481 ? _T_6887_66 : _GEN_144; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_146 = 11'h43 == _T_481 ? _T_6887_67 : _GEN_145; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_147 = 11'h44 == _T_481 ? _T_6887_68 : _GEN_146; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_148 = 11'h45 == _T_481 ? _T_6887_69 : _GEN_147; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_149 = 11'h46 == _T_481 ? _T_6887_70 : _GEN_148; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_150 = 11'h47 == _T_481 ? _T_6887_71 : _GEN_149; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_151 = 11'h48 == _T_481 ? _T_6887_72 : _GEN_150; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_152 = 11'h49 == _T_481 ? _T_6887_73 : _GEN_151; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_153 = 11'h4a == _T_481 ? _T_6887_74 : _GEN_152; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_154 = 11'h4b == _T_481 ? _T_6887_75 : _GEN_153; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_155 = 11'h4c == _T_481 ? _T_6887_76 : _GEN_154; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_156 = 11'h4d == _T_481 ? _T_6887_77 : _GEN_155; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_157 = 11'h4e == _T_481 ? _T_6887_78 : _GEN_156; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_158 = 11'h4f == _T_481 ? _T_6887_79 : _GEN_157; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_159 = 11'h50 == _T_481 ? _T_6887_80 : _GEN_158; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_160 = 11'h51 == _T_481 ? _T_6887_81 : _GEN_159; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_161 = 11'h52 == _T_481 ? _T_6887_82 : _GEN_160; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_162 = 11'h53 == _T_481 ? _T_6887_83 : _GEN_161; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_163 = 11'h54 == _T_481 ? _T_6887_84 : _GEN_162; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_164 = 11'h55 == _T_481 ? _T_6887_85 : _GEN_163; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_165 = 11'h56 == _T_481 ? _T_6887_86 : _GEN_164; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_166 = 11'h57 == _T_481 ? _T_6887_87 : _GEN_165; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_167 = 11'h58 == _T_481 ? _T_6887_88 : _GEN_166; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_168 = 11'h59 == _T_481 ? _T_6887_89 : _GEN_167; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_169 = 11'h5a == _T_481 ? _T_6887_90 : _GEN_168; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_170 = 11'h5b == _T_481 ? _T_6887_91 : _GEN_169; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_171 = 11'h5c == _T_481 ? _T_6887_92 : _GEN_170; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_172 = 11'h5d == _T_481 ? _T_6887_93 : _GEN_171; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_173 = 11'h5e == _T_481 ? _T_6887_94 : _GEN_172; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_174 = 11'h5f == _T_481 ? _T_6887_95 : _GEN_173; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_175 = 11'h60 == _T_481 ? _T_6887_96 : _GEN_174; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_176 = 11'h61 == _T_481 ? _T_6887_97 : _GEN_175; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_177 = 11'h62 == _T_481 ? _T_6887_98 : _GEN_176; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_178 = 11'h63 == _T_481 ? _T_6887_99 : _GEN_177; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_179 = 11'h64 == _T_481 ? _T_6887_100 : _GEN_178; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_180 = 11'h65 == _T_481 ? _T_6887_101 : _GEN_179; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_181 = 11'h66 == _T_481 ? _T_6887_102 : _GEN_180; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_182 = 11'h67 == _T_481 ? _T_6887_103 : _GEN_181; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_183 = 11'h68 == _T_481 ? _T_6887_104 : _GEN_182; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_184 = 11'h69 == _T_481 ? _T_6887_105 : _GEN_183; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_185 = 11'h6a == _T_481 ? _T_6887_106 : _GEN_184; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_186 = 11'h6b == _T_481 ? _T_6887_107 : _GEN_185; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_187 = 11'h6c == _T_481 ? _T_6887_108 : _GEN_186; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_188 = 11'h6d == _T_481 ? _T_6887_109 : _GEN_187; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_189 = 11'h6e == _T_481 ? _T_6887_110 : _GEN_188; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_190 = 11'h6f == _T_481 ? _T_6887_111 : _GEN_189; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_191 = 11'h70 == _T_481 ? _T_6887_112 : _GEN_190; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_192 = 11'h71 == _T_481 ? _T_6887_113 : _GEN_191; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_193 = 11'h72 == _T_481 ? _T_6887_114 : _GEN_192; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_194 = 11'h73 == _T_481 ? _T_6887_115 : _GEN_193; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_195 = 11'h74 == _T_481 ? _T_6887_116 : _GEN_194; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_196 = 11'h75 == _T_481 ? _T_6887_117 : _GEN_195; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_197 = 11'h76 == _T_481 ? _T_6887_118 : _GEN_196; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_198 = 11'h77 == _T_481 ? _T_6887_119 : _GEN_197; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_199 = 11'h78 == _T_481 ? _T_6887_120 : _GEN_198; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_200 = 11'h79 == _T_481 ? _T_6887_121 : _GEN_199; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_201 = 11'h7a == _T_481 ? _T_6887_122 : _GEN_200; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_202 = 11'h7b == _T_481 ? _T_6887_123 : _GEN_201; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_203 = 11'h7c == _T_481 ? _T_6887_124 : _GEN_202; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_204 = 11'h7d == _T_481 ? _T_6887_125 : _GEN_203; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_205 = 11'h7e == _T_481 ? _T_6887_126 : _GEN_204; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_206 = 11'h7f == _T_481 ? _T_6887_127 : _GEN_205; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_207 = 11'h80 == _T_481 ? _T_6887_128 : _GEN_206; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_208 = 11'h81 == _T_481 ? _T_6887_129 : _GEN_207; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_209 = 11'h82 == _T_481 ? _T_6887_130 : _GEN_208; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_210 = 11'h83 == _T_481 ? _T_6887_131 : _GEN_209; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_211 = 11'h84 == _T_481 ? _T_6887_132 : _GEN_210; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_212 = 11'h85 == _T_481 ? _T_6887_133 : _GEN_211; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_213 = 11'h86 == _T_481 ? _T_6887_134 : _GEN_212; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_214 = 11'h87 == _T_481 ? _T_6887_135 : _GEN_213; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_215 = 11'h88 == _T_481 ? _T_6887_136 : _GEN_214; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_216 = 11'h89 == _T_481 ? _T_6887_137 : _GEN_215; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_217 = 11'h8a == _T_481 ? _T_6887_138 : _GEN_216; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_218 = 11'h8b == _T_481 ? _T_6887_139 : _GEN_217; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_219 = 11'h8c == _T_481 ? _T_6887_140 : _GEN_218; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_220 = 11'h8d == _T_481 ? _T_6887_141 : _GEN_219; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_221 = 11'h8e == _T_481 ? _T_6887_142 : _GEN_220; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_222 = 11'h8f == _T_481 ? _T_6887_143 : _GEN_221; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_223 = 11'h90 == _T_481 ? _T_6887_144 : _GEN_222; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_224 = 11'h91 == _T_481 ? _T_6887_145 : _GEN_223; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_225 = 11'h92 == _T_481 ? _T_6887_146 : _GEN_224; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_226 = 11'h93 == _T_481 ? _T_6887_147 : _GEN_225; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_227 = 11'h94 == _T_481 ? _T_6887_148 : _GEN_226; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_228 = 11'h95 == _T_481 ? _T_6887_149 : _GEN_227; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_229 = 11'h96 == _T_481 ? _T_6887_150 : _GEN_228; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_230 = 11'h97 == _T_481 ? _T_6887_151 : _GEN_229; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_231 = 11'h98 == _T_481 ? _T_6887_152 : _GEN_230; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_232 = 11'h99 == _T_481 ? _T_6887_153 : _GEN_231; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_233 = 11'h9a == _T_481 ? _T_6887_154 : _GEN_232; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_234 = 11'h9b == _T_481 ? _T_6887_155 : _GEN_233; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_235 = 11'h9c == _T_481 ? _T_6887_156 : _GEN_234; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_236 = 11'h9d == _T_481 ? _T_6887_157 : _GEN_235; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_237 = 11'h9e == _T_481 ? _T_6887_158 : _GEN_236; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_238 = 11'h9f == _T_481 ? _T_6887_159 : _GEN_237; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_239 = 11'ha0 == _T_481 ? _T_6887_160 : _GEN_238; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_240 = 11'ha1 == _T_481 ? _T_6887_161 : _GEN_239; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_241 = 11'ha2 == _T_481 ? _T_6887_162 : _GEN_240; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_242 = 11'ha3 == _T_481 ? _T_6887_163 : _GEN_241; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_243 = 11'ha4 == _T_481 ? _T_6887_164 : _GEN_242; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_244 = 11'ha5 == _T_481 ? _T_6887_165 : _GEN_243; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_245 = 11'ha6 == _T_481 ? _T_6887_166 : _GEN_244; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_246 = 11'ha7 == _T_481 ? _T_6887_167 : _GEN_245; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_247 = 11'ha8 == _T_481 ? _T_6887_168 : _GEN_246; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_248 = 11'ha9 == _T_481 ? _T_6887_169 : _GEN_247; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_249 = 11'haa == _T_481 ? _T_6887_170 : _GEN_248; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_250 = 11'hab == _T_481 ? _T_6887_171 : _GEN_249; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_251 = 11'hac == _T_481 ? _T_6887_172 : _GEN_250; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_252 = 11'had == _T_481 ? _T_6887_173 : _GEN_251; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_253 = 11'hae == _T_481 ? _T_6887_174 : _GEN_252; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_254 = 11'haf == _T_481 ? _T_6887_175 : _GEN_253; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_255 = 11'hb0 == _T_481 ? _T_6887_176 : _GEN_254; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_256 = 11'hb1 == _T_481 ? _T_6887_177 : _GEN_255; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_257 = 11'hb2 == _T_481 ? _T_6887_178 : _GEN_256; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_258 = 11'hb3 == _T_481 ? _T_6887_179 : _GEN_257; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_259 = 11'hb4 == _T_481 ? _T_6887_180 : _GEN_258; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_260 = 11'hb5 == _T_481 ? _T_6887_181 : _GEN_259; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_261 = 11'hb6 == _T_481 ? _T_6887_182 : _GEN_260; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_262 = 11'hb7 == _T_481 ? _T_6887_183 : _GEN_261; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_263 = 11'hb8 == _T_481 ? _T_6887_184 : _GEN_262; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_264 = 11'hb9 == _T_481 ? _T_6887_185 : _GEN_263; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_265 = 11'hba == _T_481 ? _T_6887_186 : _GEN_264; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_266 = 11'hbb == _T_481 ? _T_6887_187 : _GEN_265; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_267 = 11'hbc == _T_481 ? _T_6887_188 : _GEN_266; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_268 = 11'hbd == _T_481 ? _T_6887_189 : _GEN_267; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_269 = 11'hbe == _T_481 ? _T_6887_190 : _GEN_268; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_270 = 11'hbf == _T_481 ? _T_6887_191 : _GEN_269; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_271 = 11'hc0 == _T_481 ? _T_6887_192 : _GEN_270; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_272 = 11'hc1 == _T_481 ? _T_6887_193 : _GEN_271; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_273 = 11'hc2 == _T_481 ? _T_6887_194 : _GEN_272; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_274 = 11'hc3 == _T_481 ? _T_6887_195 : _GEN_273; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_275 = 11'hc4 == _T_481 ? _T_6887_196 : _GEN_274; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_276 = 11'hc5 == _T_481 ? _T_6887_197 : _GEN_275; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_277 = 11'hc6 == _T_481 ? _T_6887_198 : _GEN_276; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_278 = 11'hc7 == _T_481 ? _T_6887_199 : _GEN_277; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_279 = 11'hc8 == _T_481 ? _T_6887_200 : _GEN_278; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_280 = 11'hc9 == _T_481 ? _T_6887_201 : _GEN_279; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_281 = 11'hca == _T_481 ? _T_6887_202 : _GEN_280; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_282 = 11'hcb == _T_481 ? _T_6887_203 : _GEN_281; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_283 = 11'hcc == _T_481 ? _T_6887_204 : _GEN_282; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_284 = 11'hcd == _T_481 ? _T_6887_205 : _GEN_283; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_285 = 11'hce == _T_481 ? _T_6887_206 : _GEN_284; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_286 = 11'hcf == _T_481 ? _T_6887_207 : _GEN_285; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_287 = 11'hd0 == _T_481 ? _T_6887_208 : _GEN_286; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_288 = 11'hd1 == _T_481 ? _T_6887_209 : _GEN_287; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_289 = 11'hd2 == _T_481 ? _T_6887_210 : _GEN_288; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_290 = 11'hd3 == _T_481 ? _T_6887_211 : _GEN_289; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_291 = 11'hd4 == _T_481 ? _T_6887_212 : _GEN_290; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_292 = 11'hd5 == _T_481 ? _T_6887_213 : _GEN_291; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_293 = 11'hd6 == _T_481 ? _T_6887_214 : _GEN_292; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_294 = 11'hd7 == _T_481 ? _T_6887_215 : _GEN_293; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_295 = 11'hd8 == _T_481 ? _T_6887_216 : _GEN_294; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_296 = 11'hd9 == _T_481 ? _T_6887_217 : _GEN_295; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_297 = 11'hda == _T_481 ? _T_6887_218 : _GEN_296; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_298 = 11'hdb == _T_481 ? _T_6887_219 : _GEN_297; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_299 = 11'hdc == _T_481 ? _T_6887_220 : _GEN_298; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_300 = 11'hdd == _T_481 ? _T_6887_221 : _GEN_299; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_301 = 11'hde == _T_481 ? _T_6887_222 : _GEN_300; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_302 = 11'hdf == _T_481 ? _T_6887_223 : _GEN_301; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_303 = 11'he0 == _T_481 ? _T_6887_224 : _GEN_302; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_304 = 11'he1 == _T_481 ? _T_6887_225 : _GEN_303; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_305 = 11'he2 == _T_481 ? _T_6887_226 : _GEN_304; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_306 = 11'he3 == _T_481 ? _T_6887_227 : _GEN_305; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_307 = 11'he4 == _T_481 ? _T_6887_228 : _GEN_306; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_308 = 11'he5 == _T_481 ? _T_6887_229 : _GEN_307; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_309 = 11'he6 == _T_481 ? _T_6887_230 : _GEN_308; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_310 = 11'he7 == _T_481 ? _T_6887_231 : _GEN_309; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_311 = 11'he8 == _T_481 ? _T_6887_232 : _GEN_310; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_312 = 11'he9 == _T_481 ? _T_6887_233 : _GEN_311; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_313 = 11'hea == _T_481 ? _T_6887_234 : _GEN_312; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_314 = 11'heb == _T_481 ? _T_6887_235 : _GEN_313; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_315 = 11'hec == _T_481 ? _T_6887_236 : _GEN_314; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_316 = 11'hed == _T_481 ? _T_6887_237 : _GEN_315; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_317 = 11'hee == _T_481 ? _T_6887_238 : _GEN_316; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_318 = 11'hef == _T_481 ? _T_6887_239 : _GEN_317; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_319 = 11'hf0 == _T_481 ? _T_6887_240 : _GEN_318; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_320 = 11'hf1 == _T_481 ? _T_6887_241 : _GEN_319; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_321 = 11'hf2 == _T_481 ? _T_6887_242 : _GEN_320; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_322 = 11'hf3 == _T_481 ? _T_6887_243 : _GEN_321; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_323 = 11'hf4 == _T_481 ? _T_6887_244 : _GEN_322; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_324 = 11'hf5 == _T_481 ? _T_6887_245 : _GEN_323; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_325 = 11'hf6 == _T_481 ? _T_6887_246 : _GEN_324; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_326 = 11'hf7 == _T_481 ? _T_6887_247 : _GEN_325; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_327 = 11'hf8 == _T_481 ? _T_6887_248 : _GEN_326; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_328 = 11'hf9 == _T_481 ? _T_6887_249 : _GEN_327; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_329 = 11'hfa == _T_481 ? _T_6887_250 : _GEN_328; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_330 = 11'hfb == _T_481 ? _T_6887_251 : _GEN_329; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_331 = 11'hfc == _T_481 ? _T_6887_252 : _GEN_330; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_332 = 11'hfd == _T_481 ? _T_6887_253 : _GEN_331; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_333 = 11'hfe == _T_481 ? _T_6887_254 : _GEN_332; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_334 = 11'hff == _T_481 ? _T_6887_255 : _GEN_333; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_335 = 11'h100 == _T_481 ? _T_6887_256 : _GEN_334; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_336 = 11'h101 == _T_481 ? _T_6887_257 : _GEN_335; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_337 = 11'h102 == _T_481 ? _T_6887_258 : _GEN_336; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_338 = 11'h103 == _T_481 ? _T_6887_259 : _GEN_337; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_339 = 11'h104 == _T_481 ? _T_6887_260 : _GEN_338; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_340 = 11'h105 == _T_481 ? _T_6887_261 : _GEN_339; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_341 = 11'h106 == _T_481 ? _T_6887_262 : _GEN_340; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_342 = 11'h107 == _T_481 ? _T_6887_263 : _GEN_341; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_343 = 11'h108 == _T_481 ? _T_6887_264 : _GEN_342; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_344 = 11'h109 == _T_481 ? _T_6887_265 : _GEN_343; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_345 = 11'h10a == _T_481 ? _T_6887_266 : _GEN_344; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_346 = 11'h10b == _T_481 ? _T_6887_267 : _GEN_345; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_347 = 11'h10c == _T_481 ? _T_6887_268 : _GEN_346; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_348 = 11'h10d == _T_481 ? _T_6887_269 : _GEN_347; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_349 = 11'h10e == _T_481 ? _T_6887_270 : _GEN_348; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_350 = 11'h10f == _T_481 ? _T_6887_271 : _GEN_349; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_351 = 11'h110 == _T_481 ? _T_6887_272 : _GEN_350; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_352 = 11'h111 == _T_481 ? _T_6887_273 : _GEN_351; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_353 = 11'h112 == _T_481 ? _T_6887_274 : _GEN_352; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_354 = 11'h113 == _T_481 ? _T_6887_275 : _GEN_353; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_355 = 11'h114 == _T_481 ? _T_6887_276 : _GEN_354; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_356 = 11'h115 == _T_481 ? _T_6887_277 : _GEN_355; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_357 = 11'h116 == _T_481 ? _T_6887_278 : _GEN_356; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_358 = 11'h117 == _T_481 ? _T_6887_279 : _GEN_357; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_359 = 11'h118 == _T_481 ? _T_6887_280 : _GEN_358; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_360 = 11'h119 == _T_481 ? _T_6887_281 : _GEN_359; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_361 = 11'h11a == _T_481 ? _T_6887_282 : _GEN_360; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_362 = 11'h11b == _T_481 ? _T_6887_283 : _GEN_361; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_363 = 11'h11c == _T_481 ? _T_6887_284 : _GEN_362; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_364 = 11'h11d == _T_481 ? _T_6887_285 : _GEN_363; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_365 = 11'h11e == _T_481 ? _T_6887_286 : _GEN_364; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_366 = 11'h11f == _T_481 ? _T_6887_287 : _GEN_365; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_367 = 11'h120 == _T_481 ? _T_6887_288 : _GEN_366; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_368 = 11'h121 == _T_481 ? _T_6887_289 : _GEN_367; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_369 = 11'h122 == _T_481 ? _T_6887_290 : _GEN_368; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_370 = 11'h123 == _T_481 ? _T_6887_291 : _GEN_369; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_371 = 11'h124 == _T_481 ? _T_6887_292 : _GEN_370; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_372 = 11'h125 == _T_481 ? _T_6887_293 : _GEN_371; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_373 = 11'h126 == _T_481 ? _T_6887_294 : _GEN_372; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_374 = 11'h127 == _T_481 ? _T_6887_295 : _GEN_373; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_375 = 11'h128 == _T_481 ? _T_6887_296 : _GEN_374; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_376 = 11'h129 == _T_481 ? _T_6887_297 : _GEN_375; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_377 = 11'h12a == _T_481 ? _T_6887_298 : _GEN_376; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_378 = 11'h12b == _T_481 ? _T_6887_299 : _GEN_377; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_379 = 11'h12c == _T_481 ? _T_6887_300 : _GEN_378; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_380 = 11'h12d == _T_481 ? _T_6887_301 : _GEN_379; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_381 = 11'h12e == _T_481 ? _T_6887_302 : _GEN_380; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_382 = 11'h12f == _T_481 ? _T_6887_303 : _GEN_381; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_383 = 11'h130 == _T_481 ? _T_6887_304 : _GEN_382; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_384 = 11'h131 == _T_481 ? _T_6887_305 : _GEN_383; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_385 = 11'h132 == _T_481 ? _T_6887_306 : _GEN_384; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_386 = 11'h133 == _T_481 ? _T_6887_307 : _GEN_385; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_387 = 11'h134 == _T_481 ? _T_6887_308 : _GEN_386; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_388 = 11'h135 == _T_481 ? _T_6887_309 : _GEN_387; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_389 = 11'h136 == _T_481 ? _T_6887_310 : _GEN_388; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_390 = 11'h137 == _T_481 ? _T_6887_311 : _GEN_389; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_391 = 11'h138 == _T_481 ? _T_6887_312 : _GEN_390; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_392 = 11'h139 == _T_481 ? _T_6887_313 : _GEN_391; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_393 = 11'h13a == _T_481 ? _T_6887_314 : _GEN_392; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_394 = 11'h13b == _T_481 ? _T_6887_315 : _GEN_393; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_395 = 11'h13c == _T_481 ? _T_6887_316 : _GEN_394; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_396 = 11'h13d == _T_481 ? _T_6887_317 : _GEN_395; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_397 = 11'h13e == _T_481 ? _T_6887_318 : _GEN_396; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_398 = 11'h13f == _T_481 ? _T_6887_319 : _GEN_397; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_399 = 11'h140 == _T_481 ? _T_6887_320 : _GEN_398; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_400 = 11'h141 == _T_481 ? _T_6887_321 : _GEN_399; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_401 = 11'h142 == _T_481 ? _T_6887_322 : _GEN_400; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_402 = 11'h143 == _T_481 ? _T_6887_323 : _GEN_401; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_403 = 11'h144 == _T_481 ? _T_6887_324 : _GEN_402; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_404 = 11'h145 == _T_481 ? _T_6887_325 : _GEN_403; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_405 = 11'h146 == _T_481 ? _T_6887_326 : _GEN_404; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_406 = 11'h147 == _T_481 ? _T_6887_327 : _GEN_405; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_407 = 11'h148 == _T_481 ? _T_6887_328 : _GEN_406; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_408 = 11'h149 == _T_481 ? _T_6887_329 : _GEN_407; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_409 = 11'h14a == _T_481 ? _T_6887_330 : _GEN_408; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_410 = 11'h14b == _T_481 ? _T_6887_331 : _GEN_409; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_411 = 11'h14c == _T_481 ? _T_6887_332 : _GEN_410; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_412 = 11'h14d == _T_481 ? _T_6887_333 : _GEN_411; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_413 = 11'h14e == _T_481 ? _T_6887_334 : _GEN_412; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_414 = 11'h14f == _T_481 ? _T_6887_335 : _GEN_413; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_415 = 11'h150 == _T_481 ? _T_6887_336 : _GEN_414; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_416 = 11'h151 == _T_481 ? _T_6887_337 : _GEN_415; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_417 = 11'h152 == _T_481 ? _T_6887_338 : _GEN_416; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_418 = 11'h153 == _T_481 ? _T_6887_339 : _GEN_417; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_419 = 11'h154 == _T_481 ? _T_6887_340 : _GEN_418; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_420 = 11'h155 == _T_481 ? _T_6887_341 : _GEN_419; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_421 = 11'h156 == _T_481 ? _T_6887_342 : _GEN_420; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_422 = 11'h157 == _T_481 ? _T_6887_343 : _GEN_421; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_423 = 11'h158 == _T_481 ? _T_6887_344 : _GEN_422; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_424 = 11'h159 == _T_481 ? _T_6887_345 : _GEN_423; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_425 = 11'h15a == _T_481 ? _T_6887_346 : _GEN_424; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_426 = 11'h15b == _T_481 ? _T_6887_347 : _GEN_425; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_427 = 11'h15c == _T_481 ? _T_6887_348 : _GEN_426; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_428 = 11'h15d == _T_481 ? _T_6887_349 : _GEN_427; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_429 = 11'h15e == _T_481 ? _T_6887_350 : _GEN_428; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_430 = 11'h15f == _T_481 ? _T_6887_351 : _GEN_429; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_431 = 11'h160 == _T_481 ? _T_6887_352 : _GEN_430; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_432 = 11'h161 == _T_481 ? _T_6887_353 : _GEN_431; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_433 = 11'h162 == _T_481 ? _T_6887_354 : _GEN_432; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_434 = 11'h163 == _T_481 ? _T_6887_355 : _GEN_433; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_435 = 11'h164 == _T_481 ? _T_6887_356 : _GEN_434; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_436 = 11'h165 == _T_481 ? _T_6887_357 : _GEN_435; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_437 = 11'h166 == _T_481 ? _T_6887_358 : _GEN_436; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_438 = 11'h167 == _T_481 ? _T_6887_359 : _GEN_437; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_439 = 11'h168 == _T_481 ? _T_6887_360 : _GEN_438; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_440 = 11'h169 == _T_481 ? _T_6887_361 : _GEN_439; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_441 = 11'h16a == _T_481 ? _T_6887_362 : _GEN_440; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_442 = 11'h16b == _T_481 ? _T_6887_363 : _GEN_441; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_443 = 11'h16c == _T_481 ? _T_6887_364 : _GEN_442; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_444 = 11'h16d == _T_481 ? _T_6887_365 : _GEN_443; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_445 = 11'h16e == _T_481 ? _T_6887_366 : _GEN_444; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_446 = 11'h16f == _T_481 ? _T_6887_367 : _GEN_445; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_447 = 11'h170 == _T_481 ? _T_6887_368 : _GEN_446; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_448 = 11'h171 == _T_481 ? _T_6887_369 : _GEN_447; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_449 = 11'h172 == _T_481 ? _T_6887_370 : _GEN_448; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_450 = 11'h173 == _T_481 ? _T_6887_371 : _GEN_449; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_451 = 11'h174 == _T_481 ? _T_6887_372 : _GEN_450; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_452 = 11'h175 == _T_481 ? _T_6887_373 : _GEN_451; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_453 = 11'h176 == _T_481 ? _T_6887_374 : _GEN_452; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_454 = 11'h177 == _T_481 ? _T_6887_375 : _GEN_453; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_455 = 11'h178 == _T_481 ? _T_6887_376 : _GEN_454; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_456 = 11'h179 == _T_481 ? _T_6887_377 : _GEN_455; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_457 = 11'h17a == _T_481 ? _T_6887_378 : _GEN_456; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_458 = 11'h17b == _T_481 ? _T_6887_379 : _GEN_457; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_459 = 11'h17c == _T_481 ? _T_6887_380 : _GEN_458; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_460 = 11'h17d == _T_481 ? _T_6887_381 : _GEN_459; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_461 = 11'h17e == _T_481 ? _T_6887_382 : _GEN_460; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_462 = 11'h17f == _T_481 ? _T_6887_383 : _GEN_461; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_463 = 11'h180 == _T_481 ? _T_6887_384 : _GEN_462; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_464 = 11'h181 == _T_481 ? _T_6887_385 : _GEN_463; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_465 = 11'h182 == _T_481 ? _T_6887_386 : _GEN_464; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_466 = 11'h183 == _T_481 ? _T_6887_387 : _GEN_465; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_467 = 11'h184 == _T_481 ? _T_6887_388 : _GEN_466; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_468 = 11'h185 == _T_481 ? _T_6887_389 : _GEN_467; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_469 = 11'h186 == _T_481 ? _T_6887_390 : _GEN_468; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_470 = 11'h187 == _T_481 ? _T_6887_391 : _GEN_469; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_471 = 11'h188 == _T_481 ? _T_6887_392 : _GEN_470; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_472 = 11'h189 == _T_481 ? _T_6887_393 : _GEN_471; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_473 = 11'h18a == _T_481 ? _T_6887_394 : _GEN_472; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_474 = 11'h18b == _T_481 ? _T_6887_395 : _GEN_473; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_475 = 11'h18c == _T_481 ? _T_6887_396 : _GEN_474; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_476 = 11'h18d == _T_481 ? _T_6887_397 : _GEN_475; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_477 = 11'h18e == _T_481 ? _T_6887_398 : _GEN_476; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_478 = 11'h18f == _T_481 ? _T_6887_399 : _GEN_477; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_479 = 11'h190 == _T_481 ? _T_6887_400 : _GEN_478; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_480 = 11'h191 == _T_481 ? _T_6887_401 : _GEN_479; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_481 = 11'h192 == _T_481 ? _T_6887_402 : _GEN_480; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_482 = 11'h193 == _T_481 ? _T_6887_403 : _GEN_481; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_483 = 11'h194 == _T_481 ? _T_6887_404 : _GEN_482; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_484 = 11'h195 == _T_481 ? _T_6887_405 : _GEN_483; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_485 = 11'h196 == _T_481 ? _T_6887_406 : _GEN_484; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_486 = 11'h197 == _T_481 ? _T_6887_407 : _GEN_485; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_487 = 11'h198 == _T_481 ? _T_6887_408 : _GEN_486; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_488 = 11'h199 == _T_481 ? _T_6887_409 : _GEN_487; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_489 = 11'h19a == _T_481 ? _T_6887_410 : _GEN_488; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_490 = 11'h19b == _T_481 ? _T_6887_411 : _GEN_489; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_491 = 11'h19c == _T_481 ? _T_6887_412 : _GEN_490; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_492 = 11'h19d == _T_481 ? _T_6887_413 : _GEN_491; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_493 = 11'h19e == _T_481 ? _T_6887_414 : _GEN_492; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_494 = 11'h19f == _T_481 ? _T_6887_415 : _GEN_493; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_495 = 11'h1a0 == _T_481 ? _T_6887_416 : _GEN_494; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_496 = 11'h1a1 == _T_481 ? _T_6887_417 : _GEN_495; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_497 = 11'h1a2 == _T_481 ? _T_6887_418 : _GEN_496; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_498 = 11'h1a3 == _T_481 ? _T_6887_419 : _GEN_497; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_499 = 11'h1a4 == _T_481 ? _T_6887_420 : _GEN_498; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_500 = 11'h1a5 == _T_481 ? _T_6887_421 : _GEN_499; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_501 = 11'h1a6 == _T_481 ? _T_6887_422 : _GEN_500; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_502 = 11'h1a7 == _T_481 ? _T_6887_423 : _GEN_501; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_503 = 11'h1a8 == _T_481 ? _T_6887_424 : _GEN_502; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_504 = 11'h1a9 == _T_481 ? _T_6887_425 : _GEN_503; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_505 = 11'h1aa == _T_481 ? _T_6887_426 : _GEN_504; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_506 = 11'h1ab == _T_481 ? _T_6887_427 : _GEN_505; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_507 = 11'h1ac == _T_481 ? _T_6887_428 : _GEN_506; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_508 = 11'h1ad == _T_481 ? _T_6887_429 : _GEN_507; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_509 = 11'h1ae == _T_481 ? _T_6887_430 : _GEN_508; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_510 = 11'h1af == _T_481 ? _T_6887_431 : _GEN_509; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_511 = 11'h1b0 == _T_481 ? _T_6887_432 : _GEN_510; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_512 = 11'h1b1 == _T_481 ? _T_6887_433 : _GEN_511; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_513 = 11'h1b2 == _T_481 ? _T_6887_434 : _GEN_512; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_514 = 11'h1b3 == _T_481 ? _T_6887_435 : _GEN_513; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_515 = 11'h1b4 == _T_481 ? _T_6887_436 : _GEN_514; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_516 = 11'h1b5 == _T_481 ? _T_6887_437 : _GEN_515; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_517 = 11'h1b6 == _T_481 ? _T_6887_438 : _GEN_516; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_518 = 11'h1b7 == _T_481 ? _T_6887_439 : _GEN_517; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_519 = 11'h1b8 == _T_481 ? _T_6887_440 : _GEN_518; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_520 = 11'h1b9 == _T_481 ? _T_6887_441 : _GEN_519; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_521 = 11'h1ba == _T_481 ? _T_6887_442 : _GEN_520; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_522 = 11'h1bb == _T_481 ? _T_6887_443 : _GEN_521; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_523 = 11'h1bc == _T_481 ? _T_6887_444 : _GEN_522; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_524 = 11'h1bd == _T_481 ? _T_6887_445 : _GEN_523; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_525 = 11'h1be == _T_481 ? _T_6887_446 : _GEN_524; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_526 = 11'h1bf == _T_481 ? _T_6887_447 : _GEN_525; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_527 = 11'h1c0 == _T_481 ? _T_6887_448 : _GEN_526; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_528 = 11'h1c1 == _T_481 ? _T_6887_449 : _GEN_527; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_529 = 11'h1c2 == _T_481 ? _T_6887_450 : _GEN_528; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_530 = 11'h1c3 == _T_481 ? _T_6887_451 : _GEN_529; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_531 = 11'h1c4 == _T_481 ? _T_6887_452 : _GEN_530; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_532 = 11'h1c5 == _T_481 ? _T_6887_453 : _GEN_531; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_533 = 11'h1c6 == _T_481 ? _T_6887_454 : _GEN_532; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_534 = 11'h1c7 == _T_481 ? _T_6887_455 : _GEN_533; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_535 = 11'h1c8 == _T_481 ? _T_6887_456 : _GEN_534; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_536 = 11'h1c9 == _T_481 ? _T_6887_457 : _GEN_535; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_537 = 11'h1ca == _T_481 ? _T_6887_458 : _GEN_536; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_538 = 11'h1cb == _T_481 ? _T_6887_459 : _GEN_537; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_539 = 11'h1cc == _T_481 ? _T_6887_460 : _GEN_538; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_540 = 11'h1cd == _T_481 ? _T_6887_461 : _GEN_539; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_541 = 11'h1ce == _T_481 ? _T_6887_462 : _GEN_540; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_542 = 11'h1cf == _T_481 ? _T_6887_463 : _GEN_541; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_543 = 11'h1d0 == _T_481 ? _T_6887_464 : _GEN_542; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_544 = 11'h1d1 == _T_481 ? _T_6887_465 : _GEN_543; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_545 = 11'h1d2 == _T_481 ? _T_6887_466 : _GEN_544; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_546 = 11'h1d3 == _T_481 ? _T_6887_467 : _GEN_545; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_547 = 11'h1d4 == _T_481 ? _T_6887_468 : _GEN_546; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_548 = 11'h1d5 == _T_481 ? _T_6887_469 : _GEN_547; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_549 = 11'h1d6 == _T_481 ? _T_6887_470 : _GEN_548; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_550 = 11'h1d7 == _T_481 ? _T_6887_471 : _GEN_549; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_551 = 11'h1d8 == _T_481 ? _T_6887_472 : _GEN_550; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_552 = 11'h1d9 == _T_481 ? _T_6887_473 : _GEN_551; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_553 = 11'h1da == _T_481 ? _T_6887_474 : _GEN_552; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_554 = 11'h1db == _T_481 ? _T_6887_475 : _GEN_553; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_555 = 11'h1dc == _T_481 ? _T_6887_476 : _GEN_554; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_556 = 11'h1dd == _T_481 ? _T_6887_477 : _GEN_555; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_557 = 11'h1de == _T_481 ? _T_6887_478 : _GEN_556; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_558 = 11'h1df == _T_481 ? _T_6887_479 : _GEN_557; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_559 = 11'h1e0 == _T_481 ? _T_6887_480 : _GEN_558; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_560 = 11'h1e1 == _T_481 ? _T_6887_481 : _GEN_559; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_561 = 11'h1e2 == _T_481 ? _T_6887_482 : _GEN_560; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_562 = 11'h1e3 == _T_481 ? _T_6887_483 : _GEN_561; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_563 = 11'h1e4 == _T_481 ? _T_6887_484 : _GEN_562; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_564 = 11'h1e5 == _T_481 ? _T_6887_485 : _GEN_563; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_565 = 11'h1e6 == _T_481 ? _T_6887_486 : _GEN_564; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_566 = 11'h1e7 == _T_481 ? _T_6887_487 : _GEN_565; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_567 = 11'h1e8 == _T_481 ? _T_6887_488 : _GEN_566; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_568 = 11'h1e9 == _T_481 ? _T_6887_489 : _GEN_567; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_569 = 11'h1ea == _T_481 ? _T_6887_490 : _GEN_568; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_570 = 11'h1eb == _T_481 ? _T_6887_491 : _GEN_569; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_571 = 11'h1ec == _T_481 ? _T_6887_492 : _GEN_570; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_572 = 11'h1ed == _T_481 ? _T_6887_493 : _GEN_571; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_573 = 11'h1ee == _T_481 ? _T_6887_494 : _GEN_572; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_574 = 11'h1ef == _T_481 ? _T_6887_495 : _GEN_573; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_575 = 11'h1f0 == _T_481 ? _T_6887_496 : _GEN_574; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_576 = 11'h1f1 == _T_481 ? _T_6887_497 : _GEN_575; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_577 = 11'h1f2 == _T_481 ? _T_6887_498 : _GEN_576; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_578 = 11'h1f3 == _T_481 ? _T_6887_499 : _GEN_577; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_579 = 11'h1f4 == _T_481 ? _T_6887_500 : _GEN_578; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_580 = 11'h1f5 == _T_481 ? _T_6887_501 : _GEN_579; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_581 = 11'h1f6 == _T_481 ? _T_6887_502 : _GEN_580; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_582 = 11'h1f7 == _T_481 ? _T_6887_503 : _GEN_581; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_583 = 11'h1f8 == _T_481 ? _T_6887_504 : _GEN_582; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_584 = 11'h1f9 == _T_481 ? _T_6887_505 : _GEN_583; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_585 = 11'h1fa == _T_481 ? _T_6887_506 : _GEN_584; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_586 = 11'h1fb == _T_481 ? _T_6887_507 : _GEN_585; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_587 = 11'h1fc == _T_481 ? _T_6887_508 : _GEN_586; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_588 = 11'h1fd == _T_481 ? _T_6887_509 : _GEN_587; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_589 = 11'h1fe == _T_481 ? _T_6887_510 : _GEN_588; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_590 = 11'h1ff == _T_481 ? _T_6887_511 : _GEN_589; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_591 = 11'h200 == _T_481 ? _T_6887_512 : _GEN_590; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_592 = 11'h201 == _T_481 ? _T_6887_513 : _GEN_591; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_593 = 11'h202 == _T_481 ? _T_6887_514 : _GEN_592; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_594 = 11'h203 == _T_481 ? _T_6887_515 : _GEN_593; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_595 = 11'h204 == _T_481 ? _T_6887_516 : _GEN_594; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_596 = 11'h205 == _T_481 ? _T_6887_517 : _GEN_595; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_597 = 11'h206 == _T_481 ? _T_6887_518 : _GEN_596; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_598 = 11'h207 == _T_481 ? _T_6887_519 : _GEN_597; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_599 = 11'h208 == _T_481 ? _T_6887_520 : _GEN_598; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_600 = 11'h209 == _T_481 ? _T_6887_521 : _GEN_599; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_601 = 11'h20a == _T_481 ? _T_6887_522 : _GEN_600; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_602 = 11'h20b == _T_481 ? _T_6887_523 : _GEN_601; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_603 = 11'h20c == _T_481 ? _T_6887_524 : _GEN_602; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_604 = 11'h20d == _T_481 ? _T_6887_525 : _GEN_603; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_605 = 11'h20e == _T_481 ? _T_6887_526 : _GEN_604; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_606 = 11'h20f == _T_481 ? _T_6887_527 : _GEN_605; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_607 = 11'h210 == _T_481 ? _T_6887_528 : _GEN_606; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_608 = 11'h211 == _T_481 ? _T_6887_529 : _GEN_607; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_609 = 11'h212 == _T_481 ? _T_6887_530 : _GEN_608; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_610 = 11'h213 == _T_481 ? _T_6887_531 : _GEN_609; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_611 = 11'h214 == _T_481 ? _T_6887_532 : _GEN_610; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_612 = 11'h215 == _T_481 ? _T_6887_533 : _GEN_611; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_613 = 11'h216 == _T_481 ? _T_6887_534 : _GEN_612; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_614 = 11'h217 == _T_481 ? _T_6887_535 : _GEN_613; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_615 = 11'h218 == _T_481 ? _T_6887_536 : _GEN_614; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_616 = 11'h219 == _T_481 ? _T_6887_537 : _GEN_615; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_617 = 11'h21a == _T_481 ? _T_6887_538 : _GEN_616; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_618 = 11'h21b == _T_481 ? _T_6887_539 : _GEN_617; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_619 = 11'h21c == _T_481 ? _T_6887_540 : _GEN_618; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_620 = 11'h21d == _T_481 ? _T_6887_541 : _GEN_619; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_621 = 11'h21e == _T_481 ? _T_6887_542 : _GEN_620; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_622 = 11'h21f == _T_481 ? _T_6887_543 : _GEN_621; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_623 = 11'h220 == _T_481 ? _T_6887_544 : _GEN_622; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_624 = 11'h221 == _T_481 ? _T_6887_545 : _GEN_623; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_625 = 11'h222 == _T_481 ? _T_6887_546 : _GEN_624; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_626 = 11'h223 == _T_481 ? _T_6887_547 : _GEN_625; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_627 = 11'h224 == _T_481 ? _T_6887_548 : _GEN_626; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_628 = 11'h225 == _T_481 ? _T_6887_549 : _GEN_627; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_629 = 11'h226 == _T_481 ? _T_6887_550 : _GEN_628; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_630 = 11'h227 == _T_481 ? _T_6887_551 : _GEN_629; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_631 = 11'h228 == _T_481 ? _T_6887_552 : _GEN_630; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_632 = 11'h229 == _T_481 ? _T_6887_553 : _GEN_631; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_633 = 11'h22a == _T_481 ? _T_6887_554 : _GEN_632; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_634 = 11'h22b == _T_481 ? _T_6887_555 : _GEN_633; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_635 = 11'h22c == _T_481 ? _T_6887_556 : _GEN_634; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_636 = 11'h22d == _T_481 ? _T_6887_557 : _GEN_635; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_637 = 11'h22e == _T_481 ? _T_6887_558 : _GEN_636; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_638 = 11'h22f == _T_481 ? _T_6887_559 : _GEN_637; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_639 = 11'h230 == _T_481 ? _T_6887_560 : _GEN_638; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_640 = 11'h231 == _T_481 ? _T_6887_561 : _GEN_639; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_641 = 11'h232 == _T_481 ? _T_6887_562 : _GEN_640; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_642 = 11'h233 == _T_481 ? _T_6887_563 : _GEN_641; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_643 = 11'h234 == _T_481 ? _T_6887_564 : _GEN_642; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_644 = 11'h235 == _T_481 ? _T_6887_565 : _GEN_643; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_645 = 11'h236 == _T_481 ? _T_6887_566 : _GEN_644; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_646 = 11'h237 == _T_481 ? _T_6887_567 : _GEN_645; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_647 = 11'h238 == _T_481 ? _T_6887_568 : _GEN_646; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_648 = 11'h239 == _T_481 ? _T_6887_569 : _GEN_647; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_649 = 11'h23a == _T_481 ? _T_6887_570 : _GEN_648; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_650 = 11'h23b == _T_481 ? _T_6887_571 : _GEN_649; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_651 = 11'h23c == _T_481 ? _T_6887_572 : _GEN_650; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_652 = 11'h23d == _T_481 ? _T_6887_573 : _GEN_651; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_653 = 11'h23e == _T_481 ? _T_6887_574 : _GEN_652; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_654 = 11'h23f == _T_481 ? _T_6887_575 : _GEN_653; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_655 = 11'h240 == _T_481 ? _T_6887_576 : _GEN_654; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_656 = 11'h241 == _T_481 ? _T_6887_577 : _GEN_655; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_657 = 11'h242 == _T_481 ? _T_6887_578 : _GEN_656; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_658 = 11'h243 == _T_481 ? _T_6887_579 : _GEN_657; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_659 = 11'h244 == _T_481 ? _T_6887_580 : _GEN_658; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_660 = 11'h245 == _T_481 ? _T_6887_581 : _GEN_659; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_661 = 11'h246 == _T_481 ? _T_6887_582 : _GEN_660; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_662 = 11'h247 == _T_481 ? _T_6887_583 : _GEN_661; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_663 = 11'h248 == _T_481 ? _T_6887_584 : _GEN_662; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_664 = 11'h249 == _T_481 ? _T_6887_585 : _GEN_663; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_665 = 11'h24a == _T_481 ? _T_6887_586 : _GEN_664; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_666 = 11'h24b == _T_481 ? _T_6887_587 : _GEN_665; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_667 = 11'h24c == _T_481 ? _T_6887_588 : _GEN_666; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_668 = 11'h24d == _T_481 ? _T_6887_589 : _GEN_667; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_669 = 11'h24e == _T_481 ? _T_6887_590 : _GEN_668; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_670 = 11'h24f == _T_481 ? _T_6887_591 : _GEN_669; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_671 = 11'h250 == _T_481 ? _T_6887_592 : _GEN_670; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_672 = 11'h251 == _T_481 ? _T_6887_593 : _GEN_671; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_673 = 11'h252 == _T_481 ? _T_6887_594 : _GEN_672; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_674 = 11'h253 == _T_481 ? _T_6887_595 : _GEN_673; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_675 = 11'h254 == _T_481 ? _T_6887_596 : _GEN_674; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_676 = 11'h255 == _T_481 ? _T_6887_597 : _GEN_675; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_677 = 11'h256 == _T_481 ? _T_6887_598 : _GEN_676; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_678 = 11'h257 == _T_481 ? _T_6887_599 : _GEN_677; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_679 = 11'h258 == _T_481 ? _T_6887_600 : _GEN_678; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_680 = 11'h259 == _T_481 ? _T_6887_601 : _GEN_679; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_681 = 11'h25a == _T_481 ? _T_6887_602 : _GEN_680; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_682 = 11'h25b == _T_481 ? _T_6887_603 : _GEN_681; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_683 = 11'h25c == _T_481 ? _T_6887_604 : _GEN_682; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_684 = 11'h25d == _T_481 ? _T_6887_605 : _GEN_683; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_685 = 11'h25e == _T_481 ? _T_6887_606 : _GEN_684; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_686 = 11'h25f == _T_481 ? _T_6887_607 : _GEN_685; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_687 = 11'h260 == _T_481 ? _T_6887_608 : _GEN_686; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_688 = 11'h261 == _T_481 ? _T_6887_609 : _GEN_687; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_689 = 11'h262 == _T_481 ? _T_6887_610 : _GEN_688; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_690 = 11'h263 == _T_481 ? _T_6887_611 : _GEN_689; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_691 = 11'h264 == _T_481 ? _T_6887_612 : _GEN_690; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_692 = 11'h265 == _T_481 ? _T_6887_613 : _GEN_691; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_693 = 11'h266 == _T_481 ? _T_6887_614 : _GEN_692; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_694 = 11'h267 == _T_481 ? _T_6887_615 : _GEN_693; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_695 = 11'h268 == _T_481 ? _T_6887_616 : _GEN_694; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_696 = 11'h269 == _T_481 ? _T_6887_617 : _GEN_695; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_697 = 11'h26a == _T_481 ? _T_6887_618 : _GEN_696; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_698 = 11'h26b == _T_481 ? _T_6887_619 : _GEN_697; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_699 = 11'h26c == _T_481 ? _T_6887_620 : _GEN_698; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_700 = 11'h26d == _T_481 ? _T_6887_621 : _GEN_699; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_701 = 11'h26e == _T_481 ? _T_6887_622 : _GEN_700; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_702 = 11'h26f == _T_481 ? _T_6887_623 : _GEN_701; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_703 = 11'h270 == _T_481 ? _T_6887_624 : _GEN_702; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_704 = 11'h271 == _T_481 ? _T_6887_625 : _GEN_703; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_705 = 11'h272 == _T_481 ? _T_6887_626 : _GEN_704; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_706 = 11'h273 == _T_481 ? _T_6887_627 : _GEN_705; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_707 = 11'h274 == _T_481 ? _T_6887_628 : _GEN_706; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_708 = 11'h275 == _T_481 ? _T_6887_629 : _GEN_707; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_709 = 11'h276 == _T_481 ? _T_6887_630 : _GEN_708; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_710 = 11'h277 == _T_481 ? _T_6887_631 : _GEN_709; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_711 = 11'h278 == _T_481 ? _T_6887_632 : _GEN_710; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_712 = 11'h279 == _T_481 ? _T_6887_633 : _GEN_711; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_713 = 11'h27a == _T_481 ? _T_6887_634 : _GEN_712; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_714 = 11'h27b == _T_481 ? _T_6887_635 : _GEN_713; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_715 = 11'h27c == _T_481 ? _T_6887_636 : _GEN_714; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_716 = 11'h27d == _T_481 ? _T_6887_637 : _GEN_715; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_717 = 11'h27e == _T_481 ? _T_6887_638 : _GEN_716; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_718 = 11'h27f == _T_481 ? _T_6887_639 : _GEN_717; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_719 = 11'h280 == _T_481 ? _T_6887_640 : _GEN_718; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_720 = 11'h281 == _T_481 ? _T_6887_641 : _GEN_719; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_721 = 11'h282 == _T_481 ? _T_6887_642 : _GEN_720; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_722 = 11'h283 == _T_481 ? _T_6887_643 : _GEN_721; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_723 = 11'h284 == _T_481 ? _T_6887_644 : _GEN_722; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_724 = 11'h285 == _T_481 ? _T_6887_645 : _GEN_723; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_725 = 11'h286 == _T_481 ? _T_6887_646 : _GEN_724; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_726 = 11'h287 == _T_481 ? _T_6887_647 : _GEN_725; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_727 = 11'h288 == _T_481 ? _T_6887_648 : _GEN_726; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_728 = 11'h289 == _T_481 ? _T_6887_649 : _GEN_727; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_729 = 11'h28a == _T_481 ? _T_6887_650 : _GEN_728; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_730 = 11'h28b == _T_481 ? _T_6887_651 : _GEN_729; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_731 = 11'h28c == _T_481 ? _T_6887_652 : _GEN_730; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_732 = 11'h28d == _T_481 ? _T_6887_653 : _GEN_731; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_733 = 11'h28e == _T_481 ? _T_6887_654 : _GEN_732; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_734 = 11'h28f == _T_481 ? _T_6887_655 : _GEN_733; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_735 = 11'h290 == _T_481 ? _T_6887_656 : _GEN_734; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_736 = 11'h291 == _T_481 ? _T_6887_657 : _GEN_735; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_737 = 11'h292 == _T_481 ? _T_6887_658 : _GEN_736; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_738 = 11'h293 == _T_481 ? _T_6887_659 : _GEN_737; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_739 = 11'h294 == _T_481 ? _T_6887_660 : _GEN_738; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_740 = 11'h295 == _T_481 ? _T_6887_661 : _GEN_739; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_741 = 11'h296 == _T_481 ? _T_6887_662 : _GEN_740; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_742 = 11'h297 == _T_481 ? _T_6887_663 : _GEN_741; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_743 = 11'h298 == _T_481 ? _T_6887_664 : _GEN_742; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_744 = 11'h299 == _T_481 ? _T_6887_665 : _GEN_743; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_745 = 11'h29a == _T_481 ? _T_6887_666 : _GEN_744; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_746 = 11'h29b == _T_481 ? _T_6887_667 : _GEN_745; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_747 = 11'h29c == _T_481 ? _T_6887_668 : _GEN_746; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_748 = 11'h29d == _T_481 ? _T_6887_669 : _GEN_747; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_749 = 11'h29e == _T_481 ? _T_6887_670 : _GEN_748; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_750 = 11'h29f == _T_481 ? _T_6887_671 : _GEN_749; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_751 = 11'h2a0 == _T_481 ? _T_6887_672 : _GEN_750; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_752 = 11'h2a1 == _T_481 ? _T_6887_673 : _GEN_751; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_753 = 11'h2a2 == _T_481 ? _T_6887_674 : _GEN_752; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_754 = 11'h2a3 == _T_481 ? _T_6887_675 : _GEN_753; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_755 = 11'h2a4 == _T_481 ? _T_6887_676 : _GEN_754; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_756 = 11'h2a5 == _T_481 ? _T_6887_677 : _GEN_755; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_757 = 11'h2a6 == _T_481 ? _T_6887_678 : _GEN_756; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_758 = 11'h2a7 == _T_481 ? _T_6887_679 : _GEN_757; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_759 = 11'h2a8 == _T_481 ? _T_6887_680 : _GEN_758; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_760 = 11'h2a9 == _T_481 ? _T_6887_681 : _GEN_759; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_761 = 11'h2aa == _T_481 ? _T_6887_682 : _GEN_760; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_762 = 11'h2ab == _T_481 ? _T_6887_683 : _GEN_761; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_763 = 11'h2ac == _T_481 ? _T_6887_684 : _GEN_762; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_764 = 11'h2ad == _T_481 ? _T_6887_685 : _GEN_763; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_765 = 11'h2ae == _T_481 ? _T_6887_686 : _GEN_764; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_766 = 11'h2af == _T_481 ? _T_6887_687 : _GEN_765; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_767 = 11'h2b0 == _T_481 ? _T_6887_688 : _GEN_766; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_768 = 11'h2b1 == _T_481 ? _T_6887_689 : _GEN_767; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_769 = 11'h2b2 == _T_481 ? _T_6887_690 : _GEN_768; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_770 = 11'h2b3 == _T_481 ? _T_6887_691 : _GEN_769; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_771 = 11'h2b4 == _T_481 ? _T_6887_692 : _GEN_770; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_772 = 11'h2b5 == _T_481 ? _T_6887_693 : _GEN_771; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_773 = 11'h2b6 == _T_481 ? _T_6887_694 : _GEN_772; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_774 = 11'h2b7 == _T_481 ? _T_6887_695 : _GEN_773; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_775 = 11'h2b8 == _T_481 ? _T_6887_696 : _GEN_774; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_776 = 11'h2b9 == _T_481 ? _T_6887_697 : _GEN_775; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_777 = 11'h2ba == _T_481 ? _T_6887_698 : _GEN_776; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_778 = 11'h2bb == _T_481 ? _T_6887_699 : _GEN_777; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_779 = 11'h2bc == _T_481 ? _T_6887_700 : _GEN_778; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_780 = 11'h2bd == _T_481 ? _T_6887_701 : _GEN_779; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_781 = 11'h2be == _T_481 ? _T_6887_702 : _GEN_780; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_782 = 11'h2bf == _T_481 ? _T_6887_703 : _GEN_781; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_783 = 11'h2c0 == _T_481 ? _T_6887_704 : _GEN_782; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_784 = 11'h2c1 == _T_481 ? _T_6887_705 : _GEN_783; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_785 = 11'h2c2 == _T_481 ? _T_6887_706 : _GEN_784; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_786 = 11'h2c3 == _T_481 ? _T_6887_707 : _GEN_785; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_787 = 11'h2c4 == _T_481 ? _T_6887_708 : _GEN_786; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_788 = 11'h2c5 == _T_481 ? _T_6887_709 : _GEN_787; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_789 = 11'h2c6 == _T_481 ? _T_6887_710 : _GEN_788; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_790 = 11'h2c7 == _T_481 ? _T_6887_711 : _GEN_789; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_791 = 11'h2c8 == _T_481 ? _T_6887_712 : _GEN_790; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_792 = 11'h2c9 == _T_481 ? _T_6887_713 : _GEN_791; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_793 = 11'h2ca == _T_481 ? _T_6887_714 : _GEN_792; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_794 = 11'h2cb == _T_481 ? _T_6887_715 : _GEN_793; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_795 = 11'h2cc == _T_481 ? _T_6887_716 : _GEN_794; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_796 = 11'h2cd == _T_481 ? _T_6887_717 : _GEN_795; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_797 = 11'h2ce == _T_481 ? _T_6887_718 : _GEN_796; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_798 = 11'h2cf == _T_481 ? _T_6887_719 : _GEN_797; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_799 = 11'h2d0 == _T_481 ? _T_6887_720 : _GEN_798; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_800 = 11'h2d1 == _T_481 ? _T_6887_721 : _GEN_799; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_801 = 11'h2d2 == _T_481 ? _T_6887_722 : _GEN_800; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_802 = 11'h2d3 == _T_481 ? _T_6887_723 : _GEN_801; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_803 = 11'h2d4 == _T_481 ? _T_6887_724 : _GEN_802; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_804 = 11'h2d5 == _T_481 ? _T_6887_725 : _GEN_803; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_805 = 11'h2d6 == _T_481 ? _T_6887_726 : _GEN_804; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_806 = 11'h2d7 == _T_481 ? _T_6887_727 : _GEN_805; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_807 = 11'h2d8 == _T_481 ? _T_6887_728 : _GEN_806; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_808 = 11'h2d9 == _T_481 ? _T_6887_729 : _GEN_807; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_809 = 11'h2da == _T_481 ? _T_6887_730 : _GEN_808; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_810 = 11'h2db == _T_481 ? _T_6887_731 : _GEN_809; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_811 = 11'h2dc == _T_481 ? _T_6887_732 : _GEN_810; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_812 = 11'h2dd == _T_481 ? _T_6887_733 : _GEN_811; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_813 = 11'h2de == _T_481 ? _T_6887_734 : _GEN_812; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_814 = 11'h2df == _T_481 ? _T_6887_735 : _GEN_813; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_815 = 11'h2e0 == _T_481 ? _T_6887_736 : _GEN_814; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_816 = 11'h2e1 == _T_481 ? _T_6887_737 : _GEN_815; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_817 = 11'h2e2 == _T_481 ? _T_6887_738 : _GEN_816; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_818 = 11'h2e3 == _T_481 ? _T_6887_739 : _GEN_817; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_819 = 11'h2e4 == _T_481 ? _T_6887_740 : _GEN_818; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_820 = 11'h2e5 == _T_481 ? _T_6887_741 : _GEN_819; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_821 = 11'h2e6 == _T_481 ? _T_6887_742 : _GEN_820; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_822 = 11'h2e7 == _T_481 ? _T_6887_743 : _GEN_821; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_823 = 11'h2e8 == _T_481 ? _T_6887_744 : _GEN_822; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_824 = 11'h2e9 == _T_481 ? _T_6887_745 : _GEN_823; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_825 = 11'h2ea == _T_481 ? _T_6887_746 : _GEN_824; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_826 = 11'h2eb == _T_481 ? _T_6887_747 : _GEN_825; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_827 = 11'h2ec == _T_481 ? _T_6887_748 : _GEN_826; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_828 = 11'h2ed == _T_481 ? _T_6887_749 : _GEN_827; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_829 = 11'h2ee == _T_481 ? _T_6887_750 : _GEN_828; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_830 = 11'h2ef == _T_481 ? _T_6887_751 : _GEN_829; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_831 = 11'h2f0 == _T_481 ? _T_6887_752 : _GEN_830; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_832 = 11'h2f1 == _T_481 ? _T_6887_753 : _GEN_831; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_833 = 11'h2f2 == _T_481 ? _T_6887_754 : _GEN_832; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_834 = 11'h2f3 == _T_481 ? _T_6887_755 : _GEN_833; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_835 = 11'h2f4 == _T_481 ? _T_6887_756 : _GEN_834; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_836 = 11'h2f5 == _T_481 ? _T_6887_757 : _GEN_835; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_837 = 11'h2f6 == _T_481 ? _T_6887_758 : _GEN_836; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_838 = 11'h2f7 == _T_481 ? _T_6887_759 : _GEN_837; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_839 = 11'h2f8 == _T_481 ? _T_6887_760 : _GEN_838; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_840 = 11'h2f9 == _T_481 ? _T_6887_761 : _GEN_839; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_841 = 11'h2fa == _T_481 ? _T_6887_762 : _GEN_840; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_842 = 11'h2fb == _T_481 ? _T_6887_763 : _GEN_841; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_843 = 11'h2fc == _T_481 ? _T_6887_764 : _GEN_842; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_844 = 11'h2fd == _T_481 ? _T_6887_765 : _GEN_843; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_845 = 11'h2fe == _T_481 ? _T_6887_766 : _GEN_844; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_846 = 11'h2ff == _T_481 ? _T_6887_767 : _GEN_845; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_847 = 11'h300 == _T_481 ? _T_6887_768 : _GEN_846; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_848 = 11'h301 == _T_481 ? _T_6887_769 : _GEN_847; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_849 = 11'h302 == _T_481 ? _T_6887_770 : _GEN_848; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_850 = 11'h303 == _T_481 ? _T_6887_771 : _GEN_849; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_851 = 11'h304 == _T_481 ? _T_6887_772 : _GEN_850; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_852 = 11'h305 == _T_481 ? _T_6887_773 : _GEN_851; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_853 = 11'h306 == _T_481 ? _T_6887_774 : _GEN_852; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_854 = 11'h307 == _T_481 ? _T_6887_775 : _GEN_853; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_855 = 11'h308 == _T_481 ? _T_6887_776 : _GEN_854; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_856 = 11'h309 == _T_481 ? _T_6887_777 : _GEN_855; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_857 = 11'h30a == _T_481 ? _T_6887_778 : _GEN_856; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_858 = 11'h30b == _T_481 ? _T_6887_779 : _GEN_857; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_859 = 11'h30c == _T_481 ? _T_6887_780 : _GEN_858; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_860 = 11'h30d == _T_481 ? _T_6887_781 : _GEN_859; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_861 = 11'h30e == _T_481 ? _T_6887_782 : _GEN_860; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_862 = 11'h30f == _T_481 ? _T_6887_783 : _GEN_861; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_863 = 11'h310 == _T_481 ? _T_6887_784 : _GEN_862; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_864 = 11'h311 == _T_481 ? _T_6887_785 : _GEN_863; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_865 = 11'h312 == _T_481 ? _T_6887_786 : _GEN_864; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_866 = 11'h313 == _T_481 ? _T_6887_787 : _GEN_865; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_867 = 11'h314 == _T_481 ? _T_6887_788 : _GEN_866; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_868 = 11'h315 == _T_481 ? _T_6887_789 : _GEN_867; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_869 = 11'h316 == _T_481 ? _T_6887_790 : _GEN_868; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_870 = 11'h317 == _T_481 ? _T_6887_791 : _GEN_869; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_871 = 11'h318 == _T_481 ? _T_6887_792 : _GEN_870; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_872 = 11'h319 == _T_481 ? _T_6887_793 : _GEN_871; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_873 = 11'h31a == _T_481 ? _T_6887_794 : _GEN_872; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_874 = 11'h31b == _T_481 ? _T_6887_795 : _GEN_873; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_875 = 11'h31c == _T_481 ? _T_6887_796 : _GEN_874; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_876 = 11'h31d == _T_481 ? _T_6887_797 : _GEN_875; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_877 = 11'h31e == _T_481 ? _T_6887_798 : _GEN_876; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_878 = 11'h31f == _T_481 ? _T_6887_799 : _GEN_877; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_879 = 11'h320 == _T_481 ? _T_6887_800 : _GEN_878; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_880 = 11'h321 == _T_481 ? _T_6887_801 : _GEN_879; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_881 = 11'h322 == _T_481 ? _T_6887_802 : _GEN_880; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_882 = 11'h323 == _T_481 ? _T_6887_803 : _GEN_881; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_883 = 11'h324 == _T_481 ? _T_6887_804 : _GEN_882; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_884 = 11'h325 == _T_481 ? _T_6887_805 : _GEN_883; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_885 = 11'h326 == _T_481 ? _T_6887_806 : _GEN_884; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_886 = 11'h327 == _T_481 ? _T_6887_807 : _GEN_885; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_887 = 11'h328 == _T_481 ? _T_6887_808 : _GEN_886; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_888 = 11'h329 == _T_481 ? _T_6887_809 : _GEN_887; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_889 = 11'h32a == _T_481 ? _T_6887_810 : _GEN_888; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_890 = 11'h32b == _T_481 ? _T_6887_811 : _GEN_889; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_891 = 11'h32c == _T_481 ? _T_6887_812 : _GEN_890; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_892 = 11'h32d == _T_481 ? _T_6887_813 : _GEN_891; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_893 = 11'h32e == _T_481 ? _T_6887_814 : _GEN_892; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_894 = 11'h32f == _T_481 ? _T_6887_815 : _GEN_893; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_895 = 11'h330 == _T_481 ? _T_6887_816 : _GEN_894; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_896 = 11'h331 == _T_481 ? _T_6887_817 : _GEN_895; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_897 = 11'h332 == _T_481 ? _T_6887_818 : _GEN_896; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_898 = 11'h333 == _T_481 ? _T_6887_819 : _GEN_897; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_899 = 11'h334 == _T_481 ? _T_6887_820 : _GEN_898; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_900 = 11'h335 == _T_481 ? _T_6887_821 : _GEN_899; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_901 = 11'h336 == _T_481 ? _T_6887_822 : _GEN_900; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_902 = 11'h337 == _T_481 ? _T_6887_823 : _GEN_901; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_903 = 11'h338 == _T_481 ? _T_6887_824 : _GEN_902; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_904 = 11'h339 == _T_481 ? _T_6887_825 : _GEN_903; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_905 = 11'h33a == _T_481 ? _T_6887_826 : _GEN_904; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_906 = 11'h33b == _T_481 ? _T_6887_827 : _GEN_905; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_907 = 11'h33c == _T_481 ? _T_6887_828 : _GEN_906; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_908 = 11'h33d == _T_481 ? _T_6887_829 : _GEN_907; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_909 = 11'h33e == _T_481 ? _T_6887_830 : _GEN_908; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_910 = 11'h33f == _T_481 ? _T_6887_831 : _GEN_909; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_911 = 11'h340 == _T_481 ? _T_6887_832 : _GEN_910; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_912 = 11'h341 == _T_481 ? _T_6887_833 : _GEN_911; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_913 = 11'h342 == _T_481 ? _T_6887_834 : _GEN_912; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_914 = 11'h343 == _T_481 ? _T_6887_835 : _GEN_913; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_915 = 11'h344 == _T_481 ? _T_6887_836 : _GEN_914; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_916 = 11'h345 == _T_481 ? _T_6887_837 : _GEN_915; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_917 = 11'h346 == _T_481 ? _T_6887_838 : _GEN_916; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_918 = 11'h347 == _T_481 ? _T_6887_839 : _GEN_917; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_919 = 11'h348 == _T_481 ? _T_6887_840 : _GEN_918; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_920 = 11'h349 == _T_481 ? _T_6887_841 : _GEN_919; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_921 = 11'h34a == _T_481 ? _T_6887_842 : _GEN_920; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_922 = 11'h34b == _T_481 ? _T_6887_843 : _GEN_921; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_923 = 11'h34c == _T_481 ? _T_6887_844 : _GEN_922; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_924 = 11'h34d == _T_481 ? _T_6887_845 : _GEN_923; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_925 = 11'h34e == _T_481 ? _T_6887_846 : _GEN_924; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_926 = 11'h34f == _T_481 ? _T_6887_847 : _GEN_925; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_927 = 11'h350 == _T_481 ? _T_6887_848 : _GEN_926; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_928 = 11'h351 == _T_481 ? _T_6887_849 : _GEN_927; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_929 = 11'h352 == _T_481 ? _T_6887_850 : _GEN_928; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_930 = 11'h353 == _T_481 ? _T_6887_851 : _GEN_929; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_931 = 11'h354 == _T_481 ? _T_6887_852 : _GEN_930; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_932 = 11'h355 == _T_481 ? _T_6887_853 : _GEN_931; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_933 = 11'h356 == _T_481 ? _T_6887_854 : _GEN_932; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_934 = 11'h357 == _T_481 ? _T_6887_855 : _GEN_933; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_935 = 11'h358 == _T_481 ? _T_6887_856 : _GEN_934; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_936 = 11'h359 == _T_481 ? _T_6887_857 : _GEN_935; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_937 = 11'h35a == _T_481 ? _T_6887_858 : _GEN_936; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_938 = 11'h35b == _T_481 ? _T_6887_859 : _GEN_937; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_939 = 11'h35c == _T_481 ? _T_6887_860 : _GEN_938; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_940 = 11'h35d == _T_481 ? _T_6887_861 : _GEN_939; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_941 = 11'h35e == _T_481 ? _T_6887_862 : _GEN_940; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_942 = 11'h35f == _T_481 ? _T_6887_863 : _GEN_941; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_943 = 11'h360 == _T_481 ? _T_6887_864 : _GEN_942; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_944 = 11'h361 == _T_481 ? _T_6887_865 : _GEN_943; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_945 = 11'h362 == _T_481 ? _T_6887_866 : _GEN_944; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_946 = 11'h363 == _T_481 ? _T_6887_867 : _GEN_945; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_947 = 11'h364 == _T_481 ? _T_6887_868 : _GEN_946; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_948 = 11'h365 == _T_481 ? _T_6887_869 : _GEN_947; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_949 = 11'h366 == _T_481 ? _T_6887_870 : _GEN_948; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_950 = 11'h367 == _T_481 ? _T_6887_871 : _GEN_949; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_951 = 11'h368 == _T_481 ? _T_6887_872 : _GEN_950; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_952 = 11'h369 == _T_481 ? _T_6887_873 : _GEN_951; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_953 = 11'h36a == _T_481 ? _T_6887_874 : _GEN_952; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_954 = 11'h36b == _T_481 ? _T_6887_875 : _GEN_953; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_955 = 11'h36c == _T_481 ? _T_6887_876 : _GEN_954; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_956 = 11'h36d == _T_481 ? _T_6887_877 : _GEN_955; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_957 = 11'h36e == _T_481 ? _T_6887_878 : _GEN_956; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_958 = 11'h36f == _T_481 ? _T_6887_879 : _GEN_957; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_959 = 11'h370 == _T_481 ? _T_6887_880 : _GEN_958; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_960 = 11'h371 == _T_481 ? _T_6887_881 : _GEN_959; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_961 = 11'h372 == _T_481 ? _T_6887_882 : _GEN_960; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_962 = 11'h373 == _T_481 ? _T_6887_883 : _GEN_961; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_963 = 11'h374 == _T_481 ? _T_6887_884 : _GEN_962; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_964 = 11'h375 == _T_481 ? _T_6887_885 : _GEN_963; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_965 = 11'h376 == _T_481 ? _T_6887_886 : _GEN_964; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_966 = 11'h377 == _T_481 ? _T_6887_887 : _GEN_965; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_967 = 11'h378 == _T_481 ? _T_6887_888 : _GEN_966; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_968 = 11'h379 == _T_481 ? _T_6887_889 : _GEN_967; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_969 = 11'h37a == _T_481 ? _T_6887_890 : _GEN_968; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_970 = 11'h37b == _T_481 ? _T_6887_891 : _GEN_969; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_971 = 11'h37c == _T_481 ? _T_6887_892 : _GEN_970; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_972 = 11'h37d == _T_481 ? _T_6887_893 : _GEN_971; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_973 = 11'h37e == _T_481 ? _T_6887_894 : _GEN_972; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_974 = 11'h37f == _T_481 ? _T_6887_895 : _GEN_973; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_975 = 11'h380 == _T_481 ? _T_6887_896 : _GEN_974; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_976 = 11'h381 == _T_481 ? _T_6887_897 : _GEN_975; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_977 = 11'h382 == _T_481 ? _T_6887_898 : _GEN_976; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_978 = 11'h383 == _T_481 ? _T_6887_899 : _GEN_977; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_979 = 11'h384 == _T_481 ? _T_6887_900 : _GEN_978; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_980 = 11'h385 == _T_481 ? _T_6887_901 : _GEN_979; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_981 = 11'h386 == _T_481 ? _T_6887_902 : _GEN_980; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_982 = 11'h387 == _T_481 ? _T_6887_903 : _GEN_981; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_983 = 11'h388 == _T_481 ? _T_6887_904 : _GEN_982; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_984 = 11'h389 == _T_481 ? _T_6887_905 : _GEN_983; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_985 = 11'h38a == _T_481 ? _T_6887_906 : _GEN_984; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_986 = 11'h38b == _T_481 ? _T_6887_907 : _GEN_985; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_987 = 11'h38c == _T_481 ? _T_6887_908 : _GEN_986; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_988 = 11'h38d == _T_481 ? _T_6887_909 : _GEN_987; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_989 = 11'h38e == _T_481 ? _T_6887_910 : _GEN_988; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_990 = 11'h38f == _T_481 ? _T_6887_911 : _GEN_989; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_991 = 11'h390 == _T_481 ? _T_6887_912 : _GEN_990; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_992 = 11'h391 == _T_481 ? _T_6887_913 : _GEN_991; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_993 = 11'h392 == _T_481 ? _T_6887_914 : _GEN_992; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_994 = 11'h393 == _T_481 ? _T_6887_915 : _GEN_993; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_995 = 11'h394 == _T_481 ? _T_6887_916 : _GEN_994; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_996 = 11'h395 == _T_481 ? _T_6887_917 : _GEN_995; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_997 = 11'h396 == _T_481 ? _T_6887_918 : _GEN_996; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_998 = 11'h397 == _T_481 ? _T_6887_919 : _GEN_997; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_999 = 11'h398 == _T_481 ? _T_6887_920 : _GEN_998; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1000 = 11'h399 == _T_481 ? _T_6887_921 : _GEN_999; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1001 = 11'h39a == _T_481 ? _T_6887_922 : _GEN_1000; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1002 = 11'h39b == _T_481 ? _T_6887_923 : _GEN_1001; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1003 = 11'h39c == _T_481 ? _T_6887_924 : _GEN_1002; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1004 = 11'h39d == _T_481 ? _T_6887_925 : _GEN_1003; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1005 = 11'h39e == _T_481 ? _T_6887_926 : _GEN_1004; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1006 = 11'h39f == _T_481 ? _T_6887_927 : _GEN_1005; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1007 = 11'h3a0 == _T_481 ? _T_6887_928 : _GEN_1006; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1008 = 11'h3a1 == _T_481 ? _T_6887_929 : _GEN_1007; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1009 = 11'h3a2 == _T_481 ? _T_6887_930 : _GEN_1008; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1010 = 11'h3a3 == _T_481 ? _T_6887_931 : _GEN_1009; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1011 = 11'h3a4 == _T_481 ? _T_6887_932 : _GEN_1010; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1012 = 11'h3a5 == _T_481 ? _T_6887_933 : _GEN_1011; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1013 = 11'h3a6 == _T_481 ? _T_6887_934 : _GEN_1012; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1014 = 11'h3a7 == _T_481 ? _T_6887_935 : _GEN_1013; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1015 = 11'h3a8 == _T_481 ? _T_6887_936 : _GEN_1014; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1016 = 11'h3a9 == _T_481 ? _T_6887_937 : _GEN_1015; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1017 = 11'h3aa == _T_481 ? _T_6887_938 : _GEN_1016; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1018 = 11'h3ab == _T_481 ? _T_6887_939 : _GEN_1017; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1019 = 11'h3ac == _T_481 ? _T_6887_940 : _GEN_1018; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1020 = 11'h3ad == _T_481 ? _T_6887_941 : _GEN_1019; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1021 = 11'h3ae == _T_481 ? _T_6887_942 : _GEN_1020; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1022 = 11'h3af == _T_481 ? _T_6887_943 : _GEN_1021; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1023 = 11'h3b0 == _T_481 ? _T_6887_944 : _GEN_1022; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1024 = 11'h3b1 == _T_481 ? _T_6887_945 : _GEN_1023; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1025 = 11'h3b2 == _T_481 ? _T_6887_946 : _GEN_1024; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1026 = 11'h3b3 == _T_481 ? _T_6887_947 : _GEN_1025; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1027 = 11'h3b4 == _T_481 ? _T_6887_948 : _GEN_1026; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1028 = 11'h3b5 == _T_481 ? _T_6887_949 : _GEN_1027; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1029 = 11'h3b6 == _T_481 ? _T_6887_950 : _GEN_1028; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1030 = 11'h3b7 == _T_481 ? _T_6887_951 : _GEN_1029; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1031 = 11'h3b8 == _T_481 ? _T_6887_952 : _GEN_1030; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1032 = 11'h3b9 == _T_481 ? _T_6887_953 : _GEN_1031; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1033 = 11'h3ba == _T_481 ? _T_6887_954 : _GEN_1032; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1034 = 11'h3bb == _T_481 ? _T_6887_955 : _GEN_1033; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1035 = 11'h3bc == _T_481 ? _T_6887_956 : _GEN_1034; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1036 = 11'h3bd == _T_481 ? _T_6887_957 : _GEN_1035; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1037 = 11'h3be == _T_481 ? _T_6887_958 : _GEN_1036; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1038 = 11'h3bf == _T_481 ? _T_6887_959 : _GEN_1037; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1039 = 11'h3c0 == _T_481 ? _T_6887_960 : _GEN_1038; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1040 = 11'h3c1 == _T_481 ? _T_6887_961 : _GEN_1039; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1041 = 11'h3c2 == _T_481 ? _T_6887_962 : _GEN_1040; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1042 = 11'h3c3 == _T_481 ? _T_6887_963 : _GEN_1041; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1043 = 11'h3c4 == _T_481 ? _T_6887_964 : _GEN_1042; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1044 = 11'h3c5 == _T_481 ? _T_6887_965 : _GEN_1043; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1045 = 11'h3c6 == _T_481 ? _T_6887_966 : _GEN_1044; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1046 = 11'h3c7 == _T_481 ? _T_6887_967 : _GEN_1045; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1047 = 11'h3c8 == _T_481 ? _T_6887_968 : _GEN_1046; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1048 = 11'h3c9 == _T_481 ? _T_6887_969 : _GEN_1047; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1049 = 11'h3ca == _T_481 ? _T_6887_970 : _GEN_1048; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1050 = 11'h3cb == _T_481 ? _T_6887_971 : _GEN_1049; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1051 = 11'h3cc == _T_481 ? _T_6887_972 : _GEN_1050; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1052 = 11'h3cd == _T_481 ? _T_6887_973 : _GEN_1051; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1053 = 11'h3ce == _T_481 ? _T_6887_974 : _GEN_1052; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1054 = 11'h3cf == _T_481 ? _T_6887_975 : _GEN_1053; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1055 = 11'h3d0 == _T_481 ? _T_6887_976 : _GEN_1054; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1056 = 11'h3d1 == _T_481 ? _T_6887_977 : _GEN_1055; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1057 = 11'h3d2 == _T_481 ? _T_6887_978 : _GEN_1056; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1058 = 11'h3d3 == _T_481 ? _T_6887_979 : _GEN_1057; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1059 = 11'h3d4 == _T_481 ? _T_6887_980 : _GEN_1058; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1060 = 11'h3d5 == _T_481 ? _T_6887_981 : _GEN_1059; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1061 = 11'h3d6 == _T_481 ? _T_6887_982 : _GEN_1060; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1062 = 11'h3d7 == _T_481 ? _T_6887_983 : _GEN_1061; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1063 = 11'h3d8 == _T_481 ? _T_6887_984 : _GEN_1062; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1064 = 11'h3d9 == _T_481 ? _T_6887_985 : _GEN_1063; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1065 = 11'h3da == _T_481 ? _T_6887_986 : _GEN_1064; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1066 = 11'h3db == _T_481 ? _T_6887_987 : _GEN_1065; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1067 = 11'h3dc == _T_481 ? _T_6887_988 : _GEN_1066; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1068 = 11'h3dd == _T_481 ? _T_6887_989 : _GEN_1067; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1069 = 11'h3de == _T_481 ? _T_6887_990 : _GEN_1068; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1070 = 11'h3df == _T_481 ? _T_6887_991 : _GEN_1069; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1071 = 11'h3e0 == _T_481 ? _T_6887_992 : _GEN_1070; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1072 = 11'h3e1 == _T_481 ? _T_6887_993 : _GEN_1071; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1073 = 11'h3e2 == _T_481 ? _T_6887_994 : _GEN_1072; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1074 = 11'h3e3 == _T_481 ? _T_6887_995 : _GEN_1073; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1075 = 11'h3e4 == _T_481 ? _T_6887_996 : _GEN_1074; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1076 = 11'h3e5 == _T_481 ? _T_6887_997 : _GEN_1075; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1077 = 11'h3e6 == _T_481 ? _T_6887_998 : _GEN_1076; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1078 = 11'h3e7 == _T_481 ? _T_6887_999 : _GEN_1077; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1079 = 11'h3e8 == _T_481 ? _T_6887_1000 : _GEN_1078; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1080 = 11'h3e9 == _T_481 ? _T_6887_1001 : _GEN_1079; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1081 = 11'h3ea == _T_481 ? _T_6887_1002 : _GEN_1080; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1082 = 11'h3eb == _T_481 ? _T_6887_1003 : _GEN_1081; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1083 = 11'h3ec == _T_481 ? _T_6887_1004 : _GEN_1082; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1084 = 11'h3ed == _T_481 ? _T_6887_1005 : _GEN_1083; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1085 = 11'h3ee == _T_481 ? _T_6887_1006 : _GEN_1084; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1086 = 11'h3ef == _T_481 ? _T_6887_1007 : _GEN_1085; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1087 = 11'h3f0 == _T_481 ? _T_6887_1008 : _GEN_1086; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1088 = 11'h3f1 == _T_481 ? _T_6887_1009 : _GEN_1087; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1089 = 11'h3f2 == _T_481 ? _T_6887_1010 : _GEN_1088; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1090 = 11'h3f3 == _T_481 ? _T_6887_1011 : _GEN_1089; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1091 = 11'h3f4 == _T_481 ? _T_6887_1012 : _GEN_1090; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1092 = 11'h3f5 == _T_481 ? _T_6887_1013 : _GEN_1091; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1093 = 11'h3f6 == _T_481 ? _T_6887_1014 : _GEN_1092; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1094 = 11'h3f7 == _T_481 ? _T_6887_1015 : _GEN_1093; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1095 = 11'h3f8 == _T_481 ? _T_6887_1016 : _GEN_1094; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1096 = 11'h3f9 == _T_481 ? _T_6887_1017 : _GEN_1095; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1097 = 11'h3fa == _T_481 ? _T_6887_1018 : _GEN_1096; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1098 = 11'h3fb == _T_481 ? _T_6887_1019 : _GEN_1097; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1099 = 11'h3fc == _T_481 ? _T_6887_1020 : _GEN_1098; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1100 = 11'h3fd == _T_481 ? _T_6887_1021 : _GEN_1099; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1101 = 11'h3fe == _T_481 ? _T_6887_1022 : _GEN_1100; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1102 = 11'h3ff == _T_481 ? _T_6887_1023 : _GEN_1101; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1103 = 11'h400 == _T_481 ? _T_6887_1024 : _GEN_1102; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1104 = 11'h401 == _T_481 ? _T_6887_1025 : _GEN_1103; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1105 = 11'h402 == _T_481 ? _T_6887_1026 : _GEN_1104; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1106 = 11'h403 == _T_481 ? _T_6887_1027 : _GEN_1105; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1107 = 11'h404 == _T_481 ? _T_6887_1028 : _GEN_1106; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1108 = 11'h405 == _T_481 ? _T_6887_1029 : _GEN_1107; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1109 = 11'h406 == _T_481 ? _T_6887_1030 : _GEN_1108; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1110 = 11'h407 == _T_481 ? _T_6887_1031 : _GEN_1109; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1111 = 11'h408 == _T_481 ? _T_6887_1032 : _GEN_1110; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1112 = 11'h409 == _T_481 ? _T_6887_1033 : _GEN_1111; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1113 = 11'h40a == _T_481 ? _T_6887_1034 : _GEN_1112; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1114 = 11'h40b == _T_481 ? _T_6887_1035 : _GEN_1113; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1115 = 11'h40c == _T_481 ? _T_6887_1036 : _GEN_1114; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1116 = 11'h40d == _T_481 ? _T_6887_1037 : _GEN_1115; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1117 = 11'h40e == _T_481 ? _T_6887_1038 : _GEN_1116; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1118 = 11'h40f == _T_481 ? _T_6887_1039 : _GEN_1117; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1119 = 11'h410 == _T_481 ? _T_6887_1040 : _GEN_1118; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1120 = 11'h411 == _T_481 ? _T_6887_1041 : _GEN_1119; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1121 = 11'h412 == _T_481 ? _T_6887_1042 : _GEN_1120; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1122 = 11'h413 == _T_481 ? _T_6887_1043 : _GEN_1121; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1123 = 11'h414 == _T_481 ? _T_6887_1044 : _GEN_1122; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1124 = 11'h415 == _T_481 ? _T_6887_1045 : _GEN_1123; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1125 = 11'h416 == _T_481 ? _T_6887_1046 : _GEN_1124; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1126 = 11'h417 == _T_481 ? _T_6887_1047 : _GEN_1125; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1127 = 11'h418 == _T_481 ? _T_6887_1048 : _GEN_1126; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1128 = 11'h419 == _T_481 ? _T_6887_1049 : _GEN_1127; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1129 = 11'h41a == _T_481 ? _T_6887_1050 : _GEN_1128; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1130 = 11'h41b == _T_481 ? _T_6887_1051 : _GEN_1129; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1131 = 11'h41c == _T_481 ? _T_6887_1052 : _GEN_1130; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1132 = 11'h41d == _T_481 ? _T_6887_1053 : _GEN_1131; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1133 = 11'h41e == _T_481 ? _T_6887_1054 : _GEN_1132; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1134 = 11'h41f == _T_481 ? _T_6887_1055 : _GEN_1133; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1135 = 11'h420 == _T_481 ? _T_6887_1056 : _GEN_1134; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1136 = 11'h421 == _T_481 ? _T_6887_1057 : _GEN_1135; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1137 = 11'h422 == _T_481 ? _T_6887_1058 : _GEN_1136; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1138 = 11'h423 == _T_481 ? _T_6887_1059 : _GEN_1137; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1139 = 11'h424 == _T_481 ? _T_6887_1060 : _GEN_1138; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1140 = 11'h425 == _T_481 ? _T_6887_1061 : _GEN_1139; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1141 = 11'h426 == _T_481 ? _T_6887_1062 : _GEN_1140; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1142 = 11'h427 == _T_481 ? _T_6887_1063 : _GEN_1141; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1143 = 11'h428 == _T_481 ? _T_6887_1064 : _GEN_1142; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1144 = 11'h429 == _T_481 ? _T_6887_1065 : _GEN_1143; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1145 = 11'h42a == _T_481 ? _T_6887_1066 : _GEN_1144; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1146 = 11'h42b == _T_481 ? _T_6887_1067 : _GEN_1145; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1147 = 11'h42c == _T_481 ? _T_6887_1068 : _GEN_1146; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1148 = 11'h42d == _T_481 ? _T_6887_1069 : _GEN_1147; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1149 = 11'h42e == _T_481 ? _T_6887_1070 : _GEN_1148; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1150 = 11'h42f == _T_481 ? _T_6887_1071 : _GEN_1149; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1151 = 11'h430 == _T_481 ? _T_6887_1072 : _GEN_1150; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1152 = 11'h431 == _T_481 ? _T_6887_1073 : _GEN_1151; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1153 = 11'h432 == _T_481 ? _T_6887_1074 : _GEN_1152; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1154 = 11'h433 == _T_481 ? _T_6887_1075 : _GEN_1153; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1155 = 11'h434 == _T_481 ? _T_6887_1076 : _GEN_1154; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1156 = 11'h435 == _T_481 ? _T_6887_1077 : _GEN_1155; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1157 = 11'h436 == _T_481 ? _T_6887_1078 : _GEN_1156; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1158 = 11'h437 == _T_481 ? _T_6887_1079 : _GEN_1157; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1159 = 11'h438 == _T_481 ? _T_6887_1080 : _GEN_1158; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1160 = 11'h439 == _T_481 ? _T_6887_1081 : _GEN_1159; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1161 = 11'h43a == _T_481 ? _T_6887_1082 : _GEN_1160; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1162 = 11'h43b == _T_481 ? _T_6887_1083 : _GEN_1161; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1163 = 11'h43c == _T_481 ? _T_6887_1084 : _GEN_1162; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1164 = 11'h43d == _T_481 ? _T_6887_1085 : _GEN_1163; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1165 = 11'h43e == _T_481 ? _T_6887_1086 : _GEN_1164; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1166 = 11'h43f == _T_481 ? _T_6887_1087 : _GEN_1165; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1167 = 11'h440 == _T_481 ? _T_6887_1088 : _GEN_1166; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1168 = 11'h441 == _T_481 ? _T_6887_1089 : _GEN_1167; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1169 = 11'h442 == _T_481 ? _T_6887_1090 : _GEN_1168; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1170 = 11'h443 == _T_481 ? _T_6887_1091 : _GEN_1169; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1171 = 11'h444 == _T_481 ? _T_6887_1092 : _GEN_1170; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1172 = 11'h445 == _T_481 ? _T_6887_1093 : _GEN_1171; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1173 = 11'h446 == _T_481 ? _T_6887_1094 : _GEN_1172; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1174 = 11'h447 == _T_481 ? _T_6887_1095 : _GEN_1173; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1175 = 11'h448 == _T_481 ? _T_6887_1096 : _GEN_1174; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1176 = 11'h449 == _T_481 ? _T_6887_1097 : _GEN_1175; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1177 = 11'h44a == _T_481 ? _T_6887_1098 : _GEN_1176; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1178 = 11'h44b == _T_481 ? _T_6887_1099 : _GEN_1177; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1179 = 11'h44c == _T_481 ? _T_6887_1100 : _GEN_1178; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1180 = 11'h44d == _T_481 ? _T_6887_1101 : _GEN_1179; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1181 = 11'h44e == _T_481 ? _T_6887_1102 : _GEN_1180; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1182 = 11'h44f == _T_481 ? _T_6887_1103 : _GEN_1181; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1183 = 11'h450 == _T_481 ? _T_6887_1104 : _GEN_1182; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1184 = 11'h451 == _T_481 ? _T_6887_1105 : _GEN_1183; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1185 = 11'h452 == _T_481 ? _T_6887_1106 : _GEN_1184; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1186 = 11'h453 == _T_481 ? _T_6887_1107 : _GEN_1185; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1187 = 11'h454 == _T_481 ? _T_6887_1108 : _GEN_1186; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1188 = 11'h455 == _T_481 ? _T_6887_1109 : _GEN_1187; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1189 = 11'h456 == _T_481 ? _T_6887_1110 : _GEN_1188; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1190 = 11'h457 == _T_481 ? _T_6887_1111 : _GEN_1189; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1191 = 11'h458 == _T_481 ? _T_6887_1112 : _GEN_1190; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1192 = 11'h459 == _T_481 ? _T_6887_1113 : _GEN_1191; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1193 = 11'h45a == _T_481 ? _T_6887_1114 : _GEN_1192; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1194 = 11'h45b == _T_481 ? _T_6887_1115 : _GEN_1193; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1195 = 11'h45c == _T_481 ? _T_6887_1116 : _GEN_1194; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1196 = 11'h45d == _T_481 ? _T_6887_1117 : _GEN_1195; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1197 = 11'h45e == _T_481 ? _T_6887_1118 : _GEN_1196; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1198 = 11'h45f == _T_481 ? _T_6887_1119 : _GEN_1197; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1199 = 11'h460 == _T_481 ? _T_6887_1120 : _GEN_1198; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1200 = 11'h461 == _T_481 ? _T_6887_1121 : _GEN_1199; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1201 = 11'h462 == _T_481 ? _T_6887_1122 : _GEN_1200; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1202 = 11'h463 == _T_481 ? _T_6887_1123 : _GEN_1201; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1203 = 11'h464 == _T_481 ? _T_6887_1124 : _GEN_1202; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1204 = 11'h465 == _T_481 ? _T_6887_1125 : _GEN_1203; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1205 = 11'h466 == _T_481 ? _T_6887_1126 : _GEN_1204; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1206 = 11'h467 == _T_481 ? _T_6887_1127 : _GEN_1205; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1207 = 11'h468 == _T_481 ? _T_6887_1128 : _GEN_1206; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1208 = 11'h469 == _T_481 ? _T_6887_1129 : _GEN_1207; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1209 = 11'h46a == _T_481 ? _T_6887_1130 : _GEN_1208; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1210 = 11'h46b == _T_481 ? _T_6887_1131 : _GEN_1209; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1211 = 11'h46c == _T_481 ? _T_6887_1132 : _GEN_1210; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1212 = 11'h46d == _T_481 ? _T_6887_1133 : _GEN_1211; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1213 = 11'h46e == _T_481 ? _T_6887_1134 : _GEN_1212; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1214 = 11'h46f == _T_481 ? _T_6887_1135 : _GEN_1213; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1215 = 11'h470 == _T_481 ? _T_6887_1136 : _GEN_1214; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1216 = 11'h471 == _T_481 ? _T_6887_1137 : _GEN_1215; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1217 = 11'h472 == _T_481 ? _T_6887_1138 : _GEN_1216; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1218 = 11'h473 == _T_481 ? _T_6887_1139 : _GEN_1217; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1219 = 11'h474 == _T_481 ? _T_6887_1140 : _GEN_1218; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1220 = 11'h475 == _T_481 ? _T_6887_1141 : _GEN_1219; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1221 = 11'h476 == _T_481 ? _T_6887_1142 : _GEN_1220; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1222 = 11'h477 == _T_481 ? _T_6887_1143 : _GEN_1221; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1223 = 11'h478 == _T_481 ? _T_6887_1144 : _GEN_1222; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1224 = 11'h479 == _T_481 ? _T_6887_1145 : _GEN_1223; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1225 = 11'h47a == _T_481 ? _T_6887_1146 : _GEN_1224; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1226 = 11'h47b == _T_481 ? _T_6887_1147 : _GEN_1225; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1227 = 11'h47c == _T_481 ? _T_6887_1148 : _GEN_1226; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1228 = 11'h47d == _T_481 ? _T_6887_1149 : _GEN_1227; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1229 = 11'h47e == _T_481 ? _T_6887_1150 : _GEN_1228; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1230 = 11'h47f == _T_481 ? _T_6887_1151 : _GEN_1229; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1231 = 11'h480 == _T_481 ? _T_6887_1152 : _GEN_1230; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1232 = 11'h481 == _T_481 ? _T_6887_1153 : _GEN_1231; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1233 = 11'h482 == _T_481 ? _T_6887_1154 : _GEN_1232; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1234 = 11'h483 == _T_481 ? _T_6887_1155 : _GEN_1233; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1235 = 11'h484 == _T_481 ? _T_6887_1156 : _GEN_1234; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1236 = 11'h485 == _T_481 ? _T_6887_1157 : _GEN_1235; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1237 = 11'h486 == _T_481 ? _T_6887_1158 : _GEN_1236; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1238 = 11'h487 == _T_481 ? _T_6887_1159 : _GEN_1237; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1239 = 11'h488 == _T_481 ? _T_6887_1160 : _GEN_1238; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1240 = 11'h489 == _T_481 ? _T_6887_1161 : _GEN_1239; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1241 = 11'h48a == _T_481 ? _T_6887_1162 : _GEN_1240; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1242 = 11'h48b == _T_481 ? _T_6887_1163 : _GEN_1241; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1243 = 11'h48c == _T_481 ? _T_6887_1164 : _GEN_1242; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1244 = 11'h48d == _T_481 ? _T_6887_1165 : _GEN_1243; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1245 = 11'h48e == _T_481 ? _T_6887_1166 : _GEN_1244; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1246 = 11'h48f == _T_481 ? _T_6887_1167 : _GEN_1245; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1247 = 11'h490 == _T_481 ? _T_6887_1168 : _GEN_1246; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1248 = 11'h491 == _T_481 ? _T_6887_1169 : _GEN_1247; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1249 = 11'h492 == _T_481 ? _T_6887_1170 : _GEN_1248; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1250 = 11'h493 == _T_481 ? _T_6887_1171 : _GEN_1249; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1251 = 11'h494 == _T_481 ? _T_6887_1172 : _GEN_1250; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1252 = 11'h495 == _T_481 ? _T_6887_1173 : _GEN_1251; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1253 = 11'h496 == _T_481 ? _T_6887_1174 : _GEN_1252; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1254 = 11'h497 == _T_481 ? _T_6887_1175 : _GEN_1253; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1255 = 11'h498 == _T_481 ? _T_6887_1176 : _GEN_1254; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1256 = 11'h499 == _T_481 ? _T_6887_1177 : _GEN_1255; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1257 = 11'h49a == _T_481 ? _T_6887_1178 : _GEN_1256; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1258 = 11'h49b == _T_481 ? _T_6887_1179 : _GEN_1257; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1259 = 11'h49c == _T_481 ? _T_6887_1180 : _GEN_1258; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1260 = 11'h49d == _T_481 ? _T_6887_1181 : _GEN_1259; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1261 = 11'h49e == _T_481 ? _T_6887_1182 : _GEN_1260; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1262 = 11'h49f == _T_481 ? _T_6887_1183 : _GEN_1261; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1263 = 11'h4a0 == _T_481 ? _T_6887_1184 : _GEN_1262; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1264 = 11'h4a1 == _T_481 ? _T_6887_1185 : _GEN_1263; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1265 = 11'h4a2 == _T_481 ? _T_6887_1186 : _GEN_1264; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1266 = 11'h4a3 == _T_481 ? _T_6887_1187 : _GEN_1265; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1267 = 11'h4a4 == _T_481 ? _T_6887_1188 : _GEN_1266; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1268 = 11'h4a5 == _T_481 ? _T_6887_1189 : _GEN_1267; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1269 = 11'h4a6 == _T_481 ? _T_6887_1190 : _GEN_1268; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1270 = 11'h4a7 == _T_481 ? _T_6887_1191 : _GEN_1269; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1271 = 11'h4a8 == _T_481 ? _T_6887_1192 : _GEN_1270; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1272 = 11'h4a9 == _T_481 ? _T_6887_1193 : _GEN_1271; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1273 = 11'h4aa == _T_481 ? _T_6887_1194 : _GEN_1272; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1274 = 11'h4ab == _T_481 ? _T_6887_1195 : _GEN_1273; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1275 = 11'h4ac == _T_481 ? _T_6887_1196 : _GEN_1274; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1276 = 11'h4ad == _T_481 ? _T_6887_1197 : _GEN_1275; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1277 = 11'h4ae == _T_481 ? _T_6887_1198 : _GEN_1276; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1278 = 11'h4af == _T_481 ? _T_6887_1199 : _GEN_1277; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1279 = 11'h4b0 == _T_481 ? _T_6887_1200 : _GEN_1278; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1280 = 11'h4b1 == _T_481 ? _T_6887_1201 : _GEN_1279; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1281 = 11'h4b2 == _T_481 ? _T_6887_1202 : _GEN_1280; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1282 = 11'h4b3 == _T_481 ? _T_6887_1203 : _GEN_1281; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1283 = 11'h4b4 == _T_481 ? _T_6887_1204 : _GEN_1282; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1284 = 11'h4b5 == _T_481 ? _T_6887_1205 : _GEN_1283; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1285 = 11'h4b6 == _T_481 ? _T_6887_1206 : _GEN_1284; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1286 = 11'h4b7 == _T_481 ? _T_6887_1207 : _GEN_1285; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1287 = 11'h4b8 == _T_481 ? _T_6887_1208 : _GEN_1286; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1288 = 11'h4b9 == _T_481 ? _T_6887_1209 : _GEN_1287; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1289 = 11'h4ba == _T_481 ? _T_6887_1210 : _GEN_1288; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1290 = 11'h4bb == _T_481 ? _T_6887_1211 : _GEN_1289; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1291 = 11'h4bc == _T_481 ? _T_6887_1212 : _GEN_1290; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1292 = 11'h4bd == _T_481 ? _T_6887_1213 : _GEN_1291; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1293 = 11'h4be == _T_481 ? _T_6887_1214 : _GEN_1292; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1294 = 11'h4bf == _T_481 ? _T_6887_1215 : _GEN_1293; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1295 = 11'h4c0 == _T_481 ? _T_6887_1216 : _GEN_1294; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1296 = 11'h4c1 == _T_481 ? _T_6887_1217 : _GEN_1295; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1297 = 11'h4c2 == _T_481 ? _T_6887_1218 : _GEN_1296; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1298 = 11'h4c3 == _T_481 ? _T_6887_1219 : _GEN_1297; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1299 = 11'h4c4 == _T_481 ? _T_6887_1220 : _GEN_1298; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1300 = 11'h4c5 == _T_481 ? _T_6887_1221 : _GEN_1299; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1301 = 11'h4c6 == _T_481 ? _T_6887_1222 : _GEN_1300; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1302 = 11'h4c7 == _T_481 ? _T_6887_1223 : _GEN_1301; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1303 = 11'h4c8 == _T_481 ? _T_6887_1224 : _GEN_1302; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1304 = 11'h4c9 == _T_481 ? _T_6887_1225 : _GEN_1303; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1305 = 11'h4ca == _T_481 ? _T_6887_1226 : _GEN_1304; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1306 = 11'h4cb == _T_481 ? _T_6887_1227 : _GEN_1305; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1307 = 11'h4cc == _T_481 ? _T_6887_1228 : _GEN_1306; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1308 = 11'h4cd == _T_481 ? _T_6887_1229 : _GEN_1307; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1309 = 11'h4ce == _T_481 ? _T_6887_1230 : _GEN_1308; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1310 = 11'h4cf == _T_481 ? _T_6887_1231 : _GEN_1309; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1311 = 11'h4d0 == _T_481 ? _T_6887_1232 : _GEN_1310; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1312 = 11'h4d1 == _T_481 ? _T_6887_1233 : _GEN_1311; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1313 = 11'h4d2 == _T_481 ? _T_6887_1234 : _GEN_1312; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1314 = 11'h4d3 == _T_481 ? _T_6887_1235 : _GEN_1313; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1315 = 11'h4d4 == _T_481 ? _T_6887_1236 : _GEN_1314; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1316 = 11'h4d5 == _T_481 ? _T_6887_1237 : _GEN_1315; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1317 = 11'h4d6 == _T_481 ? _T_6887_1238 : _GEN_1316; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1318 = 11'h4d7 == _T_481 ? _T_6887_1239 : _GEN_1317; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1319 = 11'h4d8 == _T_481 ? _T_6887_1240 : _GEN_1318; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1320 = 11'h4d9 == _T_481 ? _T_6887_1241 : _GEN_1319; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1321 = 11'h4da == _T_481 ? _T_6887_1242 : _GEN_1320; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1322 = 11'h4db == _T_481 ? _T_6887_1243 : _GEN_1321; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1323 = 11'h4dc == _T_481 ? _T_6887_1244 : _GEN_1322; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1324 = 11'h4dd == _T_481 ? _T_6887_1245 : _GEN_1323; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1325 = 11'h4de == _T_481 ? _T_6887_1246 : _GEN_1324; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1326 = 11'h4df == _T_481 ? _T_6887_1247 : _GEN_1325; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1327 = 11'h4e0 == _T_481 ? _T_6887_1248 : _GEN_1326; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1328 = 11'h4e1 == _T_481 ? _T_6887_1249 : _GEN_1327; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1329 = 11'h4e2 == _T_481 ? _T_6887_1250 : _GEN_1328; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1330 = 11'h4e3 == _T_481 ? _T_6887_1251 : _GEN_1329; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1331 = 11'h4e4 == _T_481 ? _T_6887_1252 : _GEN_1330; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1332 = 11'h4e5 == _T_481 ? _T_6887_1253 : _GEN_1331; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1333 = 11'h4e6 == _T_481 ? _T_6887_1254 : _GEN_1332; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1334 = 11'h4e7 == _T_481 ? _T_6887_1255 : _GEN_1333; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1335 = 11'h4e8 == _T_481 ? _T_6887_1256 : _GEN_1334; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1336 = 11'h4e9 == _T_481 ? _T_6887_1257 : _GEN_1335; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1337 = 11'h4ea == _T_481 ? _T_6887_1258 : _GEN_1336; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1338 = 11'h4eb == _T_481 ? _T_6887_1259 : _GEN_1337; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1339 = 11'h4ec == _T_481 ? _T_6887_1260 : _GEN_1338; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1340 = 11'h4ed == _T_481 ? _T_6887_1261 : _GEN_1339; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1341 = 11'h4ee == _T_481 ? _T_6887_1262 : _GEN_1340; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1342 = 11'h4ef == _T_481 ? _T_6887_1263 : _GEN_1341; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1343 = 11'h4f0 == _T_481 ? _T_6887_1264 : _GEN_1342; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1344 = 11'h4f1 == _T_481 ? _T_6887_1265 : _GEN_1343; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1345 = 11'h4f2 == _T_481 ? _T_6887_1266 : _GEN_1344; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1346 = 11'h4f3 == _T_481 ? _T_6887_1267 : _GEN_1345; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1347 = 11'h4f4 == _T_481 ? _T_6887_1268 : _GEN_1346; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1348 = 11'h4f5 == _T_481 ? _T_6887_1269 : _GEN_1347; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1349 = 11'h4f6 == _T_481 ? _T_6887_1270 : _GEN_1348; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1350 = 11'h4f7 == _T_481 ? _T_6887_1271 : _GEN_1349; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1351 = 11'h4f8 == _T_481 ? _T_6887_1272 : _GEN_1350; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1352 = 11'h4f9 == _T_481 ? _T_6887_1273 : _GEN_1351; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1353 = 11'h4fa == _T_481 ? _T_6887_1274 : _GEN_1352; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1354 = 11'h4fb == _T_481 ? _T_6887_1275 : _GEN_1353; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1355 = 11'h4fc == _T_481 ? _T_6887_1276 : _GEN_1354; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1356 = 11'h4fd == _T_481 ? _T_6887_1277 : _GEN_1355; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1357 = 11'h4fe == _T_481 ? _T_6887_1278 : _GEN_1356; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1358 = 11'h4ff == _T_481 ? _T_6887_1279 : _GEN_1357; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1359 = 11'h500 == _T_481 ? _T_6887_1280 : _GEN_1358; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1360 = 11'h501 == _T_481 ? _T_6887_1281 : _GEN_1359; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1361 = 11'h502 == _T_481 ? _T_6887_1282 : _GEN_1360; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1362 = 11'h503 == _T_481 ? _T_6887_1283 : _GEN_1361; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1363 = 11'h504 == _T_481 ? _T_6887_1284 : _GEN_1362; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1364 = 11'h505 == _T_481 ? _T_6887_1285 : _GEN_1363; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1365 = 11'h506 == _T_481 ? _T_6887_1286 : _GEN_1364; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1366 = 11'h507 == _T_481 ? _T_6887_1287 : _GEN_1365; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1367 = 11'h508 == _T_481 ? _T_6887_1288 : _GEN_1366; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1368 = 11'h509 == _T_481 ? _T_6887_1289 : _GEN_1367; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1369 = 11'h50a == _T_481 ? _T_6887_1290 : _GEN_1368; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1370 = 11'h50b == _T_481 ? _T_6887_1291 : _GEN_1369; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1371 = 11'h50c == _T_481 ? _T_6887_1292 : _GEN_1370; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1372 = 11'h50d == _T_481 ? _T_6887_1293 : _GEN_1371; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1373 = 11'h50e == _T_481 ? _T_6887_1294 : _GEN_1372; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1374 = 11'h50f == _T_481 ? _T_6887_1295 : _GEN_1373; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1375 = 11'h510 == _T_481 ? _T_6887_1296 : _GEN_1374; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1376 = 11'h511 == _T_481 ? _T_6887_1297 : _GEN_1375; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1377 = 11'h512 == _T_481 ? _T_6887_1298 : _GEN_1376; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1378 = 11'h513 == _T_481 ? _T_6887_1299 : _GEN_1377; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1379 = 11'h514 == _T_481 ? _T_6887_1300 : _GEN_1378; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1380 = 11'h515 == _T_481 ? _T_6887_1301 : _GEN_1379; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1381 = 11'h516 == _T_481 ? _T_6887_1302 : _GEN_1380; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1382 = 11'h517 == _T_481 ? _T_6887_1303 : _GEN_1381; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1383 = 11'h518 == _T_481 ? _T_6887_1304 : _GEN_1382; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1384 = 11'h519 == _T_481 ? _T_6887_1305 : _GEN_1383; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1385 = 11'h51a == _T_481 ? _T_6887_1306 : _GEN_1384; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1386 = 11'h51b == _T_481 ? _T_6887_1307 : _GEN_1385; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1387 = 11'h51c == _T_481 ? _T_6887_1308 : _GEN_1386; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1388 = 11'h51d == _T_481 ? _T_6887_1309 : _GEN_1387; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1389 = 11'h51e == _T_481 ? _T_6887_1310 : _GEN_1388; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1390 = 11'h51f == _T_481 ? _T_6887_1311 : _GEN_1389; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1391 = 11'h520 == _T_481 ? _T_6887_1312 : _GEN_1390; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1392 = 11'h521 == _T_481 ? _T_6887_1313 : _GEN_1391; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1393 = 11'h522 == _T_481 ? _T_6887_1314 : _GEN_1392; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1394 = 11'h523 == _T_481 ? _T_6887_1315 : _GEN_1393; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1395 = 11'h524 == _T_481 ? _T_6887_1316 : _GEN_1394; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1396 = 11'h525 == _T_481 ? _T_6887_1317 : _GEN_1395; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1397 = 11'h526 == _T_481 ? _T_6887_1318 : _GEN_1396; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1398 = 11'h527 == _T_481 ? _T_6887_1319 : _GEN_1397; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1399 = 11'h528 == _T_481 ? _T_6887_1320 : _GEN_1398; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1400 = 11'h529 == _T_481 ? _T_6887_1321 : _GEN_1399; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1401 = 11'h52a == _T_481 ? _T_6887_1322 : _GEN_1400; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1402 = 11'h52b == _T_481 ? _T_6887_1323 : _GEN_1401; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1403 = 11'h52c == _T_481 ? _T_6887_1324 : _GEN_1402; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1404 = 11'h52d == _T_481 ? _T_6887_1325 : _GEN_1403; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1405 = 11'h52e == _T_481 ? _T_6887_1326 : _GEN_1404; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1406 = 11'h52f == _T_481 ? _T_6887_1327 : _GEN_1405; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1407 = 11'h530 == _T_481 ? _T_6887_1328 : _GEN_1406; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1408 = 11'h531 == _T_481 ? _T_6887_1329 : _GEN_1407; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1409 = 11'h532 == _T_481 ? _T_6887_1330 : _GEN_1408; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1410 = 11'h533 == _T_481 ? _T_6887_1331 : _GEN_1409; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1411 = 11'h534 == _T_481 ? _T_6887_1332 : _GEN_1410; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1412 = 11'h535 == _T_481 ? _T_6887_1333 : _GEN_1411; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1413 = 11'h536 == _T_481 ? _T_6887_1334 : _GEN_1412; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1414 = 11'h537 == _T_481 ? _T_6887_1335 : _GEN_1413; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1415 = 11'h538 == _T_481 ? _T_6887_1336 : _GEN_1414; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1416 = 11'h539 == _T_481 ? _T_6887_1337 : _GEN_1415; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1417 = 11'h53a == _T_481 ? _T_6887_1338 : _GEN_1416; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1418 = 11'h53b == _T_481 ? _T_6887_1339 : _GEN_1417; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1419 = 11'h53c == _T_481 ? _T_6887_1340 : _GEN_1418; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1420 = 11'h53d == _T_481 ? _T_6887_1341 : _GEN_1419; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1421 = 11'h53e == _T_481 ? _T_6887_1342 : _GEN_1420; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1422 = 11'h53f == _T_481 ? _T_6887_1343 : _GEN_1421; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1423 = 11'h540 == _T_481 ? _T_6887_1344 : _GEN_1422; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1424 = 11'h541 == _T_481 ? _T_6887_1345 : _GEN_1423; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1425 = 11'h542 == _T_481 ? _T_6887_1346 : _GEN_1424; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1426 = 11'h543 == _T_481 ? _T_6887_1347 : _GEN_1425; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1427 = 11'h544 == _T_481 ? _T_6887_1348 : _GEN_1426; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1428 = 11'h545 == _T_481 ? _T_6887_1349 : _GEN_1427; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1429 = 11'h546 == _T_481 ? _T_6887_1350 : _GEN_1428; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1430 = 11'h547 == _T_481 ? _T_6887_1351 : _GEN_1429; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1431 = 11'h548 == _T_481 ? _T_6887_1352 : _GEN_1430; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1432 = 11'h549 == _T_481 ? _T_6887_1353 : _GEN_1431; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1433 = 11'h54a == _T_481 ? _T_6887_1354 : _GEN_1432; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1434 = 11'h54b == _T_481 ? _T_6887_1355 : _GEN_1433; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1435 = 11'h54c == _T_481 ? _T_6887_1356 : _GEN_1434; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1436 = 11'h54d == _T_481 ? _T_6887_1357 : _GEN_1435; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1437 = 11'h54e == _T_481 ? _T_6887_1358 : _GEN_1436; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1438 = 11'h54f == _T_481 ? _T_6887_1359 : _GEN_1437; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1439 = 11'h550 == _T_481 ? _T_6887_1360 : _GEN_1438; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1440 = 11'h551 == _T_481 ? _T_6887_1361 : _GEN_1439; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1441 = 11'h552 == _T_481 ? _T_6887_1362 : _GEN_1440; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1442 = 11'h553 == _T_481 ? _T_6887_1363 : _GEN_1441; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1443 = 11'h554 == _T_481 ? _T_6887_1364 : _GEN_1442; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1444 = 11'h555 == _T_481 ? _T_6887_1365 : _GEN_1443; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1445 = 11'h556 == _T_481 ? _T_6887_1366 : _GEN_1444; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1446 = 11'h557 == _T_481 ? _T_6887_1367 : _GEN_1445; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1447 = 11'h558 == _T_481 ? _T_6887_1368 : _GEN_1446; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1448 = 11'h559 == _T_481 ? _T_6887_1369 : _GEN_1447; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1449 = 11'h55a == _T_481 ? _T_6887_1370 : _GEN_1448; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1450 = 11'h55b == _T_481 ? _T_6887_1371 : _GEN_1449; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1451 = 11'h55c == _T_481 ? _T_6887_1372 : _GEN_1450; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1452 = 11'h55d == _T_481 ? _T_6887_1373 : _GEN_1451; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1453 = 11'h55e == _T_481 ? _T_6887_1374 : _GEN_1452; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1454 = 11'h55f == _T_481 ? _T_6887_1375 : _GEN_1453; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1455 = 11'h560 == _T_481 ? _T_6887_1376 : _GEN_1454; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1456 = 11'h561 == _T_481 ? _T_6887_1377 : _GEN_1455; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1457 = 11'h562 == _T_481 ? _T_6887_1378 : _GEN_1456; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1458 = 11'h563 == _T_481 ? _T_6887_1379 : _GEN_1457; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1459 = 11'h564 == _T_481 ? _T_6887_1380 : _GEN_1458; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1460 = 11'h565 == _T_481 ? _T_6887_1381 : _GEN_1459; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1461 = 11'h566 == _T_481 ? _T_6887_1382 : _GEN_1460; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1462 = 11'h567 == _T_481 ? _T_6887_1383 : _GEN_1461; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1463 = 11'h568 == _T_481 ? _T_6887_1384 : _GEN_1462; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1464 = 11'h569 == _T_481 ? _T_6887_1385 : _GEN_1463; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1465 = 11'h56a == _T_481 ? _T_6887_1386 : _GEN_1464; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1466 = 11'h56b == _T_481 ? _T_6887_1387 : _GEN_1465; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1467 = 11'h56c == _T_481 ? _T_6887_1388 : _GEN_1466; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1468 = 11'h56d == _T_481 ? _T_6887_1389 : _GEN_1467; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1469 = 11'h56e == _T_481 ? _T_6887_1390 : _GEN_1468; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1470 = 11'h56f == _T_481 ? _T_6887_1391 : _GEN_1469; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1471 = 11'h570 == _T_481 ? _T_6887_1392 : _GEN_1470; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1472 = 11'h571 == _T_481 ? _T_6887_1393 : _GEN_1471; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1473 = 11'h572 == _T_481 ? _T_6887_1394 : _GEN_1472; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1474 = 11'h573 == _T_481 ? _T_6887_1395 : _GEN_1473; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1475 = 11'h574 == _T_481 ? _T_6887_1396 : _GEN_1474; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1476 = 11'h575 == _T_481 ? _T_6887_1397 : _GEN_1475; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1477 = 11'h576 == _T_481 ? _T_6887_1398 : _GEN_1476; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1478 = 11'h577 == _T_481 ? _T_6887_1399 : _GEN_1477; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1479 = 11'h578 == _T_481 ? _T_6887_1400 : _GEN_1478; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1480 = 11'h579 == _T_481 ? _T_6887_1401 : _GEN_1479; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1481 = 11'h57a == _T_481 ? _T_6887_1402 : _GEN_1480; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1482 = 11'h57b == _T_481 ? _T_6887_1403 : _GEN_1481; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1483 = 11'h57c == _T_481 ? _T_6887_1404 : _GEN_1482; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1484 = 11'h57d == _T_481 ? _T_6887_1405 : _GEN_1483; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1485 = 11'h57e == _T_481 ? _T_6887_1406 : _GEN_1484; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1486 = 11'h57f == _T_481 ? _T_6887_1407 : _GEN_1485; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1487 = 11'h580 == _T_481 ? _T_6887_1408 : _GEN_1486; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1488 = 11'h581 == _T_481 ? _T_6887_1409 : _GEN_1487; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1489 = 11'h582 == _T_481 ? _T_6887_1410 : _GEN_1488; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1490 = 11'h583 == _T_481 ? _T_6887_1411 : _GEN_1489; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1491 = 11'h584 == _T_481 ? _T_6887_1412 : _GEN_1490; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1492 = 11'h585 == _T_481 ? _T_6887_1413 : _GEN_1491; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1493 = 11'h586 == _T_481 ? _T_6887_1414 : _GEN_1492; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1494 = 11'h587 == _T_481 ? _T_6887_1415 : _GEN_1493; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1495 = 11'h588 == _T_481 ? _T_6887_1416 : _GEN_1494; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1496 = 11'h589 == _T_481 ? _T_6887_1417 : _GEN_1495; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1497 = 11'h58a == _T_481 ? _T_6887_1418 : _GEN_1496; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1498 = 11'h58b == _T_481 ? _T_6887_1419 : _GEN_1497; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1499 = 11'h58c == _T_481 ? _T_6887_1420 : _GEN_1498; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1500 = 11'h58d == _T_481 ? _T_6887_1421 : _GEN_1499; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1501 = 11'h58e == _T_481 ? _T_6887_1422 : _GEN_1500; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1502 = 11'h58f == _T_481 ? _T_6887_1423 : _GEN_1501; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1503 = 11'h590 == _T_481 ? _T_6887_1424 : _GEN_1502; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1504 = 11'h591 == _T_481 ? _T_6887_1425 : _GEN_1503; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1505 = 11'h592 == _T_481 ? _T_6887_1426 : _GEN_1504; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1506 = 11'h593 == _T_481 ? _T_6887_1427 : _GEN_1505; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1507 = 11'h594 == _T_481 ? _T_6887_1428 : _GEN_1506; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1508 = 11'h595 == _T_481 ? _T_6887_1429 : _GEN_1507; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1509 = 11'h596 == _T_481 ? _T_6887_1430 : _GEN_1508; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1510 = 11'h597 == _T_481 ? _T_6887_1431 : _GEN_1509; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1511 = 11'h598 == _T_481 ? _T_6887_1432 : _GEN_1510; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1512 = 11'h599 == _T_481 ? _T_6887_1433 : _GEN_1511; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1513 = 11'h59a == _T_481 ? _T_6887_1434 : _GEN_1512; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1514 = 11'h59b == _T_481 ? _T_6887_1435 : _GEN_1513; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1515 = 11'h59c == _T_481 ? _T_6887_1436 : _GEN_1514; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1516 = 11'h59d == _T_481 ? _T_6887_1437 : _GEN_1515; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1517 = 11'h59e == _T_481 ? _T_6887_1438 : _GEN_1516; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1518 = 11'h59f == _T_481 ? _T_6887_1439 : _GEN_1517; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1519 = 11'h5a0 == _T_481 ? _T_6887_1440 : _GEN_1518; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1520 = 11'h5a1 == _T_481 ? _T_6887_1441 : _GEN_1519; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1521 = 11'h5a2 == _T_481 ? _T_6887_1442 : _GEN_1520; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1522 = 11'h5a3 == _T_481 ? _T_6887_1443 : _GEN_1521; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1523 = 11'h5a4 == _T_481 ? _T_6887_1444 : _GEN_1522; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1524 = 11'h5a5 == _T_481 ? _T_6887_1445 : _GEN_1523; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1525 = 11'h5a6 == _T_481 ? _T_6887_1446 : _GEN_1524; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1526 = 11'h5a7 == _T_481 ? _T_6887_1447 : _GEN_1525; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1527 = 11'h5a8 == _T_481 ? _T_6887_1448 : _GEN_1526; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1528 = 11'h5a9 == _T_481 ? _T_6887_1449 : _GEN_1527; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1529 = 11'h5aa == _T_481 ? _T_6887_1450 : _GEN_1528; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1530 = 11'h5ab == _T_481 ? _T_6887_1451 : _GEN_1529; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1531 = 11'h5ac == _T_481 ? _T_6887_1452 : _GEN_1530; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1532 = 11'h5ad == _T_481 ? _T_6887_1453 : _GEN_1531; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1533 = 11'h5ae == _T_481 ? _T_6887_1454 : _GEN_1532; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1534 = 11'h5af == _T_481 ? _T_6887_1455 : _GEN_1533; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1535 = 11'h5b0 == _T_481 ? _T_6887_1456 : _GEN_1534; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1536 = 11'h5b1 == _T_481 ? _T_6887_1457 : _GEN_1535; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1537 = 11'h5b2 == _T_481 ? _T_6887_1458 : _GEN_1536; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1538 = 11'h5b3 == _T_481 ? _T_6887_1459 : _GEN_1537; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1539 = 11'h5b4 == _T_481 ? _T_6887_1460 : _GEN_1538; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1540 = 11'h5b5 == _T_481 ? _T_6887_1461 : _GEN_1539; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1541 = 11'h5b6 == _T_481 ? _T_6887_1462 : _GEN_1540; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1542 = 11'h5b7 == _T_481 ? _T_6887_1463 : _GEN_1541; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1543 = 11'h5b8 == _T_481 ? _T_6887_1464 : _GEN_1542; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1544 = 11'h5b9 == _T_481 ? _T_6887_1465 : _GEN_1543; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1545 = 11'h5ba == _T_481 ? _T_6887_1466 : _GEN_1544; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1546 = 11'h5bb == _T_481 ? _T_6887_1467 : _GEN_1545; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1547 = 11'h5bc == _T_481 ? _T_6887_1468 : _GEN_1546; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1548 = 11'h5bd == _T_481 ? _T_6887_1469 : _GEN_1547; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1549 = 11'h5be == _T_481 ? _T_6887_1470 : _GEN_1548; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1550 = 11'h5bf == _T_481 ? _T_6887_1471 : _GEN_1549; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1551 = 11'h5c0 == _T_481 ? _T_6887_1472 : _GEN_1550; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1552 = 11'h5c1 == _T_481 ? _T_6887_1473 : _GEN_1551; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1553 = 11'h5c2 == _T_481 ? _T_6887_1474 : _GEN_1552; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1554 = 11'h5c3 == _T_481 ? _T_6887_1475 : _GEN_1553; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1555 = 11'h5c4 == _T_481 ? _T_6887_1476 : _GEN_1554; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1556 = 11'h5c5 == _T_481 ? _T_6887_1477 : _GEN_1555; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1557 = 11'h5c6 == _T_481 ? _T_6887_1478 : _GEN_1556; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1558 = 11'h5c7 == _T_481 ? _T_6887_1479 : _GEN_1557; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1559 = 11'h5c8 == _T_481 ? _T_6887_1480 : _GEN_1558; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1560 = 11'h5c9 == _T_481 ? _T_6887_1481 : _GEN_1559; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1561 = 11'h5ca == _T_481 ? _T_6887_1482 : _GEN_1560; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1562 = 11'h5cb == _T_481 ? _T_6887_1483 : _GEN_1561; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1563 = 11'h5cc == _T_481 ? _T_6887_1484 : _GEN_1562; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1564 = 11'h5cd == _T_481 ? _T_6887_1485 : _GEN_1563; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1565 = 11'h5ce == _T_481 ? _T_6887_1486 : _GEN_1564; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1566 = 11'h5cf == _T_481 ? _T_6887_1487 : _GEN_1565; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1567 = 11'h5d0 == _T_481 ? _T_6887_1488 : _GEN_1566; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1568 = 11'h5d1 == _T_481 ? _T_6887_1489 : _GEN_1567; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1569 = 11'h5d2 == _T_481 ? _T_6887_1490 : _GEN_1568; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1570 = 11'h5d3 == _T_481 ? _T_6887_1491 : _GEN_1569; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1571 = 11'h5d4 == _T_481 ? _T_6887_1492 : _GEN_1570; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1572 = 11'h5d5 == _T_481 ? _T_6887_1493 : _GEN_1571; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1573 = 11'h5d6 == _T_481 ? _T_6887_1494 : _GEN_1572; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1574 = 11'h5d7 == _T_481 ? _T_6887_1495 : _GEN_1573; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1575 = 11'h5d8 == _T_481 ? _T_6887_1496 : _GEN_1574; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1576 = 11'h5d9 == _T_481 ? _T_6887_1497 : _GEN_1575; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1577 = 11'h5da == _T_481 ? _T_6887_1498 : _GEN_1576; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1578 = 11'h5db == _T_481 ? _T_6887_1499 : _GEN_1577; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1579 = 11'h5dc == _T_481 ? _T_6887_1500 : _GEN_1578; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1580 = 11'h5dd == _T_481 ? _T_6887_1501 : _GEN_1579; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1581 = 11'h5de == _T_481 ? _T_6887_1502 : _GEN_1580; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1582 = 11'h5df == _T_481 ? _T_6887_1503 : _GEN_1581; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1583 = 11'h5e0 == _T_481 ? _T_6887_1504 : _GEN_1582; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1584 = 11'h5e1 == _T_481 ? _T_6887_1505 : _GEN_1583; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1585 = 11'h5e2 == _T_481 ? _T_6887_1506 : _GEN_1584; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1586 = 11'h5e3 == _T_481 ? _T_6887_1507 : _GEN_1585; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1587 = 11'h5e4 == _T_481 ? _T_6887_1508 : _GEN_1586; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1588 = 11'h5e5 == _T_481 ? _T_6887_1509 : _GEN_1587; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1589 = 11'h5e6 == _T_481 ? _T_6887_1510 : _GEN_1588; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1590 = 11'h5e7 == _T_481 ? _T_6887_1511 : _GEN_1589; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1591 = 11'h5e8 == _T_481 ? _T_6887_1512 : _GEN_1590; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1592 = 11'h5e9 == _T_481 ? _T_6887_1513 : _GEN_1591; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1593 = 11'h5ea == _T_481 ? _T_6887_1514 : _GEN_1592; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1594 = 11'h5eb == _T_481 ? _T_6887_1515 : _GEN_1593; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1595 = 11'h5ec == _T_481 ? _T_6887_1516 : _GEN_1594; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1596 = 11'h5ed == _T_481 ? _T_6887_1517 : _GEN_1595; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1597 = 11'h5ee == _T_481 ? _T_6887_1518 : _GEN_1596; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1598 = 11'h5ef == _T_481 ? _T_6887_1519 : _GEN_1597; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1599 = 11'h5f0 == _T_481 ? _T_6887_1520 : _GEN_1598; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1600 = 11'h5f1 == _T_481 ? _T_6887_1521 : _GEN_1599; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1601 = 11'h5f2 == _T_481 ? _T_6887_1522 : _GEN_1600; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1602 = 11'h5f3 == _T_481 ? _T_6887_1523 : _GEN_1601; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1603 = 11'h5f4 == _T_481 ? _T_6887_1524 : _GEN_1602; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1604 = 11'h5f5 == _T_481 ? _T_6887_1525 : _GEN_1603; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1605 = 11'h5f6 == _T_481 ? _T_6887_1526 : _GEN_1604; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1606 = 11'h5f7 == _T_481 ? _T_6887_1527 : _GEN_1605; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1607 = 11'h5f8 == _T_481 ? _T_6887_1528 : _GEN_1606; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1608 = 11'h5f9 == _T_481 ? _T_6887_1529 : _GEN_1607; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1609 = 11'h5fa == _T_481 ? _T_6887_1530 : _GEN_1608; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1610 = 11'h5fb == _T_481 ? _T_6887_1531 : _GEN_1609; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1611 = 11'h5fc == _T_481 ? _T_6887_1532 : _GEN_1610; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1612 = 11'h5fd == _T_481 ? _T_6887_1533 : _GEN_1611; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1613 = 11'h5fe == _T_481 ? _T_6887_1534 : _GEN_1612; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1614 = 11'h5ff == _T_481 ? _T_6887_1535 : _GEN_1613; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1615 = 11'h600 == _T_481 ? _T_6887_1536 : _GEN_1614; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1616 = 11'h601 == _T_481 ? _T_6887_1537 : _GEN_1615; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1617 = 11'h602 == _T_481 ? _T_6887_1538 : _GEN_1616; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1618 = 11'h603 == _T_481 ? _T_6887_1539 : _GEN_1617; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1619 = 11'h604 == _T_481 ? _T_6887_1540 : _GEN_1618; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1620 = 11'h605 == _T_481 ? _T_6887_1541 : _GEN_1619; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1621 = 11'h606 == _T_481 ? _T_6887_1542 : _GEN_1620; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1622 = 11'h607 == _T_481 ? _T_6887_1543 : _GEN_1621; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1623 = 11'h608 == _T_481 ? _T_6887_1544 : _GEN_1622; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1624 = 11'h609 == _T_481 ? _T_6887_1545 : _GEN_1623; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1625 = 11'h60a == _T_481 ? _T_6887_1546 : _GEN_1624; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1626 = 11'h60b == _T_481 ? _T_6887_1547 : _GEN_1625; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1627 = 11'h60c == _T_481 ? _T_6887_1548 : _GEN_1626; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1628 = 11'h60d == _T_481 ? _T_6887_1549 : _GEN_1627; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1629 = 11'h60e == _T_481 ? _T_6887_1550 : _GEN_1628; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1630 = 11'h60f == _T_481 ? _T_6887_1551 : _GEN_1629; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1631 = 11'h610 == _T_481 ? _T_6887_1552 : _GEN_1630; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1632 = 11'h611 == _T_481 ? _T_6887_1553 : _GEN_1631; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1633 = 11'h612 == _T_481 ? _T_6887_1554 : _GEN_1632; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1634 = 11'h613 == _T_481 ? _T_6887_1555 : _GEN_1633; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1635 = 11'h614 == _T_481 ? _T_6887_1556 : _GEN_1634; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1636 = 11'h615 == _T_481 ? _T_6887_1557 : _GEN_1635; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1637 = 11'h616 == _T_481 ? _T_6887_1558 : _GEN_1636; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1638 = 11'h617 == _T_481 ? _T_6887_1559 : _GEN_1637; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1639 = 11'h618 == _T_481 ? _T_6887_1560 : _GEN_1638; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1640 = 11'h619 == _T_481 ? _T_6887_1561 : _GEN_1639; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1641 = 11'h61a == _T_481 ? _T_6887_1562 : _GEN_1640; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1642 = 11'h61b == _T_481 ? _T_6887_1563 : _GEN_1641; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1643 = 11'h61c == _T_481 ? _T_6887_1564 : _GEN_1642; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1644 = 11'h61d == _T_481 ? _T_6887_1565 : _GEN_1643; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1645 = 11'h61e == _T_481 ? _T_6887_1566 : _GEN_1644; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1646 = 11'h61f == _T_481 ? _T_6887_1567 : _GEN_1645; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1647 = 11'h620 == _T_481 ? _T_6887_1568 : _GEN_1646; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1648 = 11'h621 == _T_481 ? _T_6887_1569 : _GEN_1647; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1649 = 11'h622 == _T_481 ? _T_6887_1570 : _GEN_1648; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1650 = 11'h623 == _T_481 ? _T_6887_1571 : _GEN_1649; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1651 = 11'h624 == _T_481 ? _T_6887_1572 : _GEN_1650; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1652 = 11'h625 == _T_481 ? _T_6887_1573 : _GEN_1651; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1653 = 11'h626 == _T_481 ? _T_6887_1574 : _GEN_1652; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1654 = 11'h627 == _T_481 ? _T_6887_1575 : _GEN_1653; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1655 = 11'h628 == _T_481 ? _T_6887_1576 : _GEN_1654; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1656 = 11'h629 == _T_481 ? _T_6887_1577 : _GEN_1655; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1657 = 11'h62a == _T_481 ? _T_6887_1578 : _GEN_1656; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1658 = 11'h62b == _T_481 ? _T_6887_1579 : _GEN_1657; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1659 = 11'h62c == _T_481 ? _T_6887_1580 : _GEN_1658; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1660 = 11'h62d == _T_481 ? _T_6887_1581 : _GEN_1659; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1661 = 11'h62e == _T_481 ? _T_6887_1582 : _GEN_1660; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1662 = 11'h62f == _T_481 ? _T_6887_1583 : _GEN_1661; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1663 = 11'h630 == _T_481 ? _T_6887_1584 : _GEN_1662; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1664 = 11'h631 == _T_481 ? _T_6887_1585 : _GEN_1663; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1665 = 11'h632 == _T_481 ? _T_6887_1586 : _GEN_1664; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1666 = 11'h633 == _T_481 ? _T_6887_1587 : _GEN_1665; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1667 = 11'h634 == _T_481 ? _T_6887_1588 : _GEN_1666; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1668 = 11'h635 == _T_481 ? _T_6887_1589 : _GEN_1667; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1669 = 11'h636 == _T_481 ? _T_6887_1590 : _GEN_1668; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1670 = 11'h637 == _T_481 ? _T_6887_1591 : _GEN_1669; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1671 = 11'h638 == _T_481 ? _T_6887_1592 : _GEN_1670; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1672 = 11'h639 == _T_481 ? _T_6887_1593 : _GEN_1671; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1673 = 11'h63a == _T_481 ? _T_6887_1594 : _GEN_1672; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1674 = 11'h63b == _T_481 ? _T_6887_1595 : _GEN_1673; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1675 = 11'h63c == _T_481 ? _T_6887_1596 : _GEN_1674; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1676 = 11'h63d == _T_481 ? _T_6887_1597 : _GEN_1675; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1677 = 11'h63e == _T_481 ? _T_6887_1598 : _GEN_1676; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1678 = 11'h63f == _T_481 ? _T_6887_1599 : _GEN_1677; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1679 = 11'h640 == _T_481 ? _T_6887_1600 : _GEN_1678; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1680 = 11'h641 == _T_481 ? _T_6887_1601 : _GEN_1679; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1681 = 11'h642 == _T_481 ? _T_6887_1602 : _GEN_1680; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1682 = 11'h643 == _T_481 ? _T_6887_1603 : _GEN_1681; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1683 = 11'h644 == _T_481 ? _T_6887_1604 : _GEN_1682; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1684 = 11'h645 == _T_481 ? _T_6887_1605 : _GEN_1683; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1685 = 11'h646 == _T_481 ? _T_6887_1606 : _GEN_1684; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1686 = 11'h647 == _T_481 ? _T_6887_1607 : _GEN_1685; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1687 = 11'h648 == _T_481 ? _T_6887_1608 : _GEN_1686; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1688 = 11'h649 == _T_481 ? _T_6887_1609 : _GEN_1687; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1689 = 11'h64a == _T_481 ? _T_6887_1610 : _GEN_1688; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1690 = 11'h64b == _T_481 ? _T_6887_1611 : _GEN_1689; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1691 = 11'h64c == _T_481 ? _T_6887_1612 : _GEN_1690; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1692 = 11'h64d == _T_481 ? _T_6887_1613 : _GEN_1691; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1693 = 11'h64e == _T_481 ? _T_6887_1614 : _GEN_1692; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1694 = 11'h64f == _T_481 ? _T_6887_1615 : _GEN_1693; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1695 = 11'h650 == _T_481 ? _T_6887_1616 : _GEN_1694; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1696 = 11'h651 == _T_481 ? _T_6887_1617 : _GEN_1695; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1697 = 11'h652 == _T_481 ? _T_6887_1618 : _GEN_1696; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1698 = 11'h653 == _T_481 ? _T_6887_1619 : _GEN_1697; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1699 = 11'h654 == _T_481 ? _T_6887_1620 : _GEN_1698; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1700 = 11'h655 == _T_481 ? _T_6887_1621 : _GEN_1699; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1701 = 11'h656 == _T_481 ? _T_6887_1622 : _GEN_1700; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1702 = 11'h657 == _T_481 ? _T_6887_1623 : _GEN_1701; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1703 = 11'h658 == _T_481 ? _T_6887_1624 : _GEN_1702; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1704 = 11'h659 == _T_481 ? _T_6887_1625 : _GEN_1703; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1705 = 11'h65a == _T_481 ? _T_6887_1626 : _GEN_1704; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1706 = 11'h65b == _T_481 ? _T_6887_1627 : _GEN_1705; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1707 = 11'h65c == _T_481 ? _T_6887_1628 : _GEN_1706; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1708 = 11'h65d == _T_481 ? _T_6887_1629 : _GEN_1707; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1709 = 11'h65e == _T_481 ? _T_6887_1630 : _GEN_1708; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1710 = 11'h65f == _T_481 ? _T_6887_1631 : _GEN_1709; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1711 = 11'h660 == _T_481 ? _T_6887_1632 : _GEN_1710; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1712 = 11'h661 == _T_481 ? _T_6887_1633 : _GEN_1711; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1713 = 11'h662 == _T_481 ? _T_6887_1634 : _GEN_1712; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1714 = 11'h663 == _T_481 ? _T_6887_1635 : _GEN_1713; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1715 = 11'h664 == _T_481 ? _T_6887_1636 : _GEN_1714; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1716 = 11'h665 == _T_481 ? _T_6887_1637 : _GEN_1715; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1717 = 11'h666 == _T_481 ? _T_6887_1638 : _GEN_1716; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1718 = 11'h667 == _T_481 ? _T_6887_1639 : _GEN_1717; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1719 = 11'h668 == _T_481 ? _T_6887_1640 : _GEN_1718; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1720 = 11'h669 == _T_481 ? _T_6887_1641 : _GEN_1719; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1721 = 11'h66a == _T_481 ? _T_6887_1642 : _GEN_1720; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1722 = 11'h66b == _T_481 ? _T_6887_1643 : _GEN_1721; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1723 = 11'h66c == _T_481 ? _T_6887_1644 : _GEN_1722; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1724 = 11'h66d == _T_481 ? _T_6887_1645 : _GEN_1723; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1725 = 11'h66e == _T_481 ? _T_6887_1646 : _GEN_1724; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1726 = 11'h66f == _T_481 ? _T_6887_1647 : _GEN_1725; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1727 = 11'h670 == _T_481 ? _T_6887_1648 : _GEN_1726; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1728 = 11'h671 == _T_481 ? _T_6887_1649 : _GEN_1727; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1729 = 11'h672 == _T_481 ? _T_6887_1650 : _GEN_1728; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1730 = 11'h673 == _T_481 ? _T_6887_1651 : _GEN_1729; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1731 = 11'h674 == _T_481 ? _T_6887_1652 : _GEN_1730; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1732 = 11'h675 == _T_481 ? _T_6887_1653 : _GEN_1731; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1733 = 11'h676 == _T_481 ? _T_6887_1654 : _GEN_1732; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1734 = 11'h677 == _T_481 ? _T_6887_1655 : _GEN_1733; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1735 = 11'h678 == _T_481 ? _T_6887_1656 : _GEN_1734; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1736 = 11'h679 == _T_481 ? _T_6887_1657 : _GEN_1735; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1737 = 11'h67a == _T_481 ? _T_6887_1658 : _GEN_1736; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1738 = 11'h67b == _T_481 ? _T_6887_1659 : _GEN_1737; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1739 = 11'h67c == _T_481 ? _T_6887_1660 : _GEN_1738; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1740 = 11'h67d == _T_481 ? _T_6887_1661 : _GEN_1739; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1741 = 11'h67e == _T_481 ? _T_6887_1662 : _GEN_1740; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1742 = 11'h67f == _T_481 ? _T_6887_1663 : _GEN_1741; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1743 = 11'h680 == _T_481 ? _T_6887_1664 : _GEN_1742; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1744 = 11'h681 == _T_481 ? _T_6887_1665 : _GEN_1743; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1745 = 11'h682 == _T_481 ? _T_6887_1666 : _GEN_1744; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1746 = 11'h683 == _T_481 ? _T_6887_1667 : _GEN_1745; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1747 = 11'h684 == _T_481 ? _T_6887_1668 : _GEN_1746; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1748 = 11'h685 == _T_481 ? _T_6887_1669 : _GEN_1747; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1749 = 11'h686 == _T_481 ? _T_6887_1670 : _GEN_1748; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1750 = 11'h687 == _T_481 ? _T_6887_1671 : _GEN_1749; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1751 = 11'h688 == _T_481 ? _T_6887_1672 : _GEN_1750; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1752 = 11'h689 == _T_481 ? _T_6887_1673 : _GEN_1751; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1753 = 11'h68a == _T_481 ? _T_6887_1674 : _GEN_1752; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1754 = 11'h68b == _T_481 ? _T_6887_1675 : _GEN_1753; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1755 = 11'h68c == _T_481 ? _T_6887_1676 : _GEN_1754; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1756 = 11'h68d == _T_481 ? _T_6887_1677 : _GEN_1755; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1757 = 11'h68e == _T_481 ? _T_6887_1678 : _GEN_1756; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1758 = 11'h68f == _T_481 ? _T_6887_1679 : _GEN_1757; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1759 = 11'h690 == _T_481 ? _T_6887_1680 : _GEN_1758; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1760 = 11'h691 == _T_481 ? _T_6887_1681 : _GEN_1759; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1761 = 11'h692 == _T_481 ? _T_6887_1682 : _GEN_1760; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1762 = 11'h693 == _T_481 ? _T_6887_1683 : _GEN_1761; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1763 = 11'h694 == _T_481 ? _T_6887_1684 : _GEN_1762; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1764 = 11'h695 == _T_481 ? _T_6887_1685 : _GEN_1763; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1765 = 11'h696 == _T_481 ? _T_6887_1686 : _GEN_1764; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1766 = 11'h697 == _T_481 ? _T_6887_1687 : _GEN_1765; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1767 = 11'h698 == _T_481 ? _T_6887_1688 : _GEN_1766; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1768 = 11'h699 == _T_481 ? _T_6887_1689 : _GEN_1767; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1769 = 11'h69a == _T_481 ? _T_6887_1690 : _GEN_1768; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1770 = 11'h69b == _T_481 ? _T_6887_1691 : _GEN_1769; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1771 = 11'h69c == _T_481 ? _T_6887_1692 : _GEN_1770; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1772 = 11'h69d == _T_481 ? _T_6887_1693 : _GEN_1771; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1773 = 11'h69e == _T_481 ? _T_6887_1694 : _GEN_1772; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1774 = 11'h69f == _T_481 ? _T_6887_1695 : _GEN_1773; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1775 = 11'h6a0 == _T_481 ? _T_6887_1696 : _GEN_1774; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1776 = 11'h6a1 == _T_481 ? _T_6887_1697 : _GEN_1775; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1777 = 11'h6a2 == _T_481 ? _T_6887_1698 : _GEN_1776; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1778 = 11'h6a3 == _T_481 ? _T_6887_1699 : _GEN_1777; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1779 = 11'h6a4 == _T_481 ? _T_6887_1700 : _GEN_1778; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1780 = 11'h6a5 == _T_481 ? _T_6887_1701 : _GEN_1779; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1781 = 11'h6a6 == _T_481 ? _T_6887_1702 : _GEN_1780; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1782 = 11'h6a7 == _T_481 ? _T_6887_1703 : _GEN_1781; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1783 = 11'h6a8 == _T_481 ? _T_6887_1704 : _GEN_1782; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1784 = 11'h6a9 == _T_481 ? _T_6887_1705 : _GEN_1783; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1785 = 11'h6aa == _T_481 ? _T_6887_1706 : _GEN_1784; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1786 = 11'h6ab == _T_481 ? _T_6887_1707 : _GEN_1785; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1787 = 11'h6ac == _T_481 ? _T_6887_1708 : _GEN_1786; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1788 = 11'h6ad == _T_481 ? _T_6887_1709 : _GEN_1787; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1789 = 11'h6ae == _T_481 ? _T_6887_1710 : _GEN_1788; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1790 = 11'h6af == _T_481 ? _T_6887_1711 : _GEN_1789; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1791 = 11'h6b0 == _T_481 ? _T_6887_1712 : _GEN_1790; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1792 = 11'h6b1 == _T_481 ? _T_6887_1713 : _GEN_1791; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1793 = 11'h6b2 == _T_481 ? _T_6887_1714 : _GEN_1792; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1794 = 11'h6b3 == _T_481 ? _T_6887_1715 : _GEN_1793; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1795 = 11'h6b4 == _T_481 ? _T_6887_1716 : _GEN_1794; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1796 = 11'h6b5 == _T_481 ? _T_6887_1717 : _GEN_1795; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1797 = 11'h6b6 == _T_481 ? _T_6887_1718 : _GEN_1796; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1798 = 11'h6b7 == _T_481 ? _T_6887_1719 : _GEN_1797; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1799 = 11'h6b8 == _T_481 ? _T_6887_1720 : _GEN_1798; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1800 = 11'h6b9 == _T_481 ? _T_6887_1721 : _GEN_1799; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1801 = 11'h6ba == _T_481 ? _T_6887_1722 : _GEN_1800; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1802 = 11'h6bb == _T_481 ? _T_6887_1723 : _GEN_1801; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1803 = 11'h6bc == _T_481 ? _T_6887_1724 : _GEN_1802; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1804 = 11'h6bd == _T_481 ? _T_6887_1725 : _GEN_1803; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1805 = 11'h6be == _T_481 ? _T_6887_1726 : _GEN_1804; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1806 = 11'h6bf == _T_481 ? _T_6887_1727 : _GEN_1805; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1807 = 11'h6c0 == _T_481 ? _T_6887_1728 : _GEN_1806; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1808 = 11'h6c1 == _T_481 ? _T_6887_1729 : _GEN_1807; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1809 = 11'h6c2 == _T_481 ? _T_6887_1730 : _GEN_1808; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1810 = 11'h6c3 == _T_481 ? _T_6887_1731 : _GEN_1809; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1811 = 11'h6c4 == _T_481 ? _T_6887_1732 : _GEN_1810; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1812 = 11'h6c5 == _T_481 ? _T_6887_1733 : _GEN_1811; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1813 = 11'h6c6 == _T_481 ? _T_6887_1734 : _GEN_1812; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1814 = 11'h6c7 == _T_481 ? _T_6887_1735 : _GEN_1813; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1815 = 11'h6c8 == _T_481 ? _T_6887_1736 : _GEN_1814; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1816 = 11'h6c9 == _T_481 ? _T_6887_1737 : _GEN_1815; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1817 = 11'h6ca == _T_481 ? _T_6887_1738 : _GEN_1816; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1818 = 11'h6cb == _T_481 ? _T_6887_1739 : _GEN_1817; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1819 = 11'h6cc == _T_481 ? _T_6887_1740 : _GEN_1818; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1820 = 11'h6cd == _T_481 ? _T_6887_1741 : _GEN_1819; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1821 = 11'h6ce == _T_481 ? _T_6887_1742 : _GEN_1820; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1822 = 11'h6cf == _T_481 ? _T_6887_1743 : _GEN_1821; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1823 = 11'h6d0 == _T_481 ? _T_6887_1744 : _GEN_1822; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1824 = 11'h6d1 == _T_481 ? _T_6887_1745 : _GEN_1823; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1825 = 11'h6d2 == _T_481 ? _T_6887_1746 : _GEN_1824; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1826 = 11'h6d3 == _T_481 ? _T_6887_1747 : _GEN_1825; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1827 = 11'h6d4 == _T_481 ? _T_6887_1748 : _GEN_1826; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1828 = 11'h6d5 == _T_481 ? _T_6887_1749 : _GEN_1827; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1829 = 11'h6d6 == _T_481 ? _T_6887_1750 : _GEN_1828; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1830 = 11'h6d7 == _T_481 ? _T_6887_1751 : _GEN_1829; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1831 = 11'h6d8 == _T_481 ? _T_6887_1752 : _GEN_1830; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1832 = 11'h6d9 == _T_481 ? _T_6887_1753 : _GEN_1831; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1833 = 11'h6da == _T_481 ? _T_6887_1754 : _GEN_1832; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1834 = 11'h6db == _T_481 ? _T_6887_1755 : _GEN_1833; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1835 = 11'h6dc == _T_481 ? _T_6887_1756 : _GEN_1834; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1836 = 11'h6dd == _T_481 ? _T_6887_1757 : _GEN_1835; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1837 = 11'h6de == _T_481 ? _T_6887_1758 : _GEN_1836; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1838 = 11'h6df == _T_481 ? _T_6887_1759 : _GEN_1837; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1839 = 11'h6e0 == _T_481 ? _T_6887_1760 : _GEN_1838; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1840 = 11'h6e1 == _T_481 ? _T_6887_1761 : _GEN_1839; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1841 = 11'h6e2 == _T_481 ? _T_6887_1762 : _GEN_1840; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1842 = 11'h6e3 == _T_481 ? _T_6887_1763 : _GEN_1841; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1843 = 11'h6e4 == _T_481 ? _T_6887_1764 : _GEN_1842; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1844 = 11'h6e5 == _T_481 ? _T_6887_1765 : _GEN_1843; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1845 = 11'h6e6 == _T_481 ? _T_6887_1766 : _GEN_1844; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1846 = 11'h6e7 == _T_481 ? _T_6887_1767 : _GEN_1845; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1847 = 11'h6e8 == _T_481 ? _T_6887_1768 : _GEN_1846; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1848 = 11'h6e9 == _T_481 ? _T_6887_1769 : _GEN_1847; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1849 = 11'h6ea == _T_481 ? _T_6887_1770 : _GEN_1848; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1850 = 11'h6eb == _T_481 ? _T_6887_1771 : _GEN_1849; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1851 = 11'h6ec == _T_481 ? _T_6887_1772 : _GEN_1850; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1852 = 11'h6ed == _T_481 ? _T_6887_1773 : _GEN_1851; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1853 = 11'h6ee == _T_481 ? _T_6887_1774 : _GEN_1852; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1854 = 11'h6ef == _T_481 ? _T_6887_1775 : _GEN_1853; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1855 = 11'h6f0 == _T_481 ? _T_6887_1776 : _GEN_1854; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1856 = 11'h6f1 == _T_481 ? _T_6887_1777 : _GEN_1855; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1857 = 11'h6f2 == _T_481 ? _T_6887_1778 : _GEN_1856; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1858 = 11'h6f3 == _T_481 ? _T_6887_1779 : _GEN_1857; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1859 = 11'h6f4 == _T_481 ? _T_6887_1780 : _GEN_1858; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1860 = 11'h6f5 == _T_481 ? _T_6887_1781 : _GEN_1859; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1861 = 11'h6f6 == _T_481 ? _T_6887_1782 : _GEN_1860; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1862 = 11'h6f7 == _T_481 ? _T_6887_1783 : _GEN_1861; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1863 = 11'h6f8 == _T_481 ? _T_6887_1784 : _GEN_1862; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1864 = 11'h6f9 == _T_481 ? _T_6887_1785 : _GEN_1863; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1865 = 11'h6fa == _T_481 ? _T_6887_1786 : _GEN_1864; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1866 = 11'h6fb == _T_481 ? _T_6887_1787 : _GEN_1865; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1867 = 11'h6fc == _T_481 ? _T_6887_1788 : _GEN_1866; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1868 = 11'h6fd == _T_481 ? _T_6887_1789 : _GEN_1867; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1869 = 11'h6fe == _T_481 ? _T_6887_1790 : _GEN_1868; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1870 = 11'h6ff == _T_481 ? _T_6887_1791 : _GEN_1869; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1871 = 11'h700 == _T_481 ? _T_6887_1792 : _GEN_1870; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1872 = 11'h701 == _T_481 ? _T_6887_1793 : _GEN_1871; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1873 = 11'h702 == _T_481 ? _T_6887_1794 : _GEN_1872; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1874 = 11'h703 == _T_481 ? _T_6887_1795 : _GEN_1873; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1875 = 11'h704 == _T_481 ? _T_6887_1796 : _GEN_1874; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1876 = 11'h705 == _T_481 ? _T_6887_1797 : _GEN_1875; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1877 = 11'h706 == _T_481 ? _T_6887_1798 : _GEN_1876; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1878 = 11'h707 == _T_481 ? _T_6887_1799 : _GEN_1877; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1879 = 11'h708 == _T_481 ? _T_6887_1800 : _GEN_1878; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1880 = 11'h709 == _T_481 ? _T_6887_1801 : _GEN_1879; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1881 = 11'h70a == _T_481 ? _T_6887_1802 : _GEN_1880; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1882 = 11'h70b == _T_481 ? _T_6887_1803 : _GEN_1881; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1883 = 11'h70c == _T_481 ? _T_6887_1804 : _GEN_1882; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1884 = 11'h70d == _T_481 ? _T_6887_1805 : _GEN_1883; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1885 = 11'h70e == _T_481 ? _T_6887_1806 : _GEN_1884; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1886 = 11'h70f == _T_481 ? _T_6887_1807 : _GEN_1885; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1887 = 11'h710 == _T_481 ? _T_6887_1808 : _GEN_1886; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1888 = 11'h711 == _T_481 ? _T_6887_1809 : _GEN_1887; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1889 = 11'h712 == _T_481 ? _T_6887_1810 : _GEN_1888; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1890 = 11'h713 == _T_481 ? _T_6887_1811 : _GEN_1889; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1891 = 11'h714 == _T_481 ? _T_6887_1812 : _GEN_1890; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1892 = 11'h715 == _T_481 ? _T_6887_1813 : _GEN_1891; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1893 = 11'h716 == _T_481 ? _T_6887_1814 : _GEN_1892; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1894 = 11'h717 == _T_481 ? _T_6887_1815 : _GEN_1893; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1895 = 11'h718 == _T_481 ? _T_6887_1816 : _GEN_1894; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1896 = 11'h719 == _T_481 ? _T_6887_1817 : _GEN_1895; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1897 = 11'h71a == _T_481 ? _T_6887_1818 : _GEN_1896; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1898 = 11'h71b == _T_481 ? _T_6887_1819 : _GEN_1897; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1899 = 11'h71c == _T_481 ? _T_6887_1820 : _GEN_1898; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1900 = 11'h71d == _T_481 ? _T_6887_1821 : _GEN_1899; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1901 = 11'h71e == _T_481 ? _T_6887_1822 : _GEN_1900; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1902 = 11'h71f == _T_481 ? _T_6887_1823 : _GEN_1901; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1903 = 11'h720 == _T_481 ? _T_6887_1824 : _GEN_1902; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1904 = 11'h721 == _T_481 ? _T_6887_1825 : _GEN_1903; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1905 = 11'h722 == _T_481 ? _T_6887_1826 : _GEN_1904; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1906 = 11'h723 == _T_481 ? _T_6887_1827 : _GEN_1905; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1907 = 11'h724 == _T_481 ? _T_6887_1828 : _GEN_1906; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1908 = 11'h725 == _T_481 ? _T_6887_1829 : _GEN_1907; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1909 = 11'h726 == _T_481 ? _T_6887_1830 : _GEN_1908; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1910 = 11'h727 == _T_481 ? _T_6887_1831 : _GEN_1909; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1911 = 11'h728 == _T_481 ? _T_6887_1832 : _GEN_1910; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1912 = 11'h729 == _T_481 ? _T_6887_1833 : _GEN_1911; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1913 = 11'h72a == _T_481 ? _T_6887_1834 : _GEN_1912; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1914 = 11'h72b == _T_481 ? _T_6887_1835 : _GEN_1913; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1915 = 11'h72c == _T_481 ? _T_6887_1836 : _GEN_1914; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1916 = 11'h72d == _T_481 ? _T_6887_1837 : _GEN_1915; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1917 = 11'h72e == _T_481 ? _T_6887_1838 : _GEN_1916; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1918 = 11'h72f == _T_481 ? _T_6887_1839 : _GEN_1917; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1919 = 11'h730 == _T_481 ? _T_6887_1840 : _GEN_1918; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1920 = 11'h731 == _T_481 ? _T_6887_1841 : _GEN_1919; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1921 = 11'h732 == _T_481 ? _T_6887_1842 : _GEN_1920; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1922 = 11'h733 == _T_481 ? _T_6887_1843 : _GEN_1921; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1923 = 11'h734 == _T_481 ? _T_6887_1844 : _GEN_1922; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1924 = 11'h735 == _T_481 ? _T_6887_1845 : _GEN_1923; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1925 = 11'h736 == _T_481 ? _T_6887_1846 : _GEN_1924; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1926 = 11'h737 == _T_481 ? _T_6887_1847 : _GEN_1925; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1927 = 11'h738 == _T_481 ? _T_6887_1848 : _GEN_1926; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1928 = 11'h739 == _T_481 ? _T_6887_1849 : _GEN_1927; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1929 = 11'h73a == _T_481 ? _T_6887_1850 : _GEN_1928; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1930 = 11'h73b == _T_481 ? _T_6887_1851 : _GEN_1929; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1931 = 11'h73c == _T_481 ? _T_6887_1852 : _GEN_1930; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1932 = 11'h73d == _T_481 ? _T_6887_1853 : _GEN_1931; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1933 = 11'h73e == _T_481 ? _T_6887_1854 : _GEN_1932; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1934 = 11'h73f == _T_481 ? _T_6887_1855 : _GEN_1933; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1935 = 11'h740 == _T_481 ? _T_6887_1856 : _GEN_1934; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1936 = 11'h741 == _T_481 ? _T_6887_1857 : _GEN_1935; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1937 = 11'h742 == _T_481 ? _T_6887_1858 : _GEN_1936; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1938 = 11'h743 == _T_481 ? _T_6887_1859 : _GEN_1937; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1939 = 11'h744 == _T_481 ? _T_6887_1860 : _GEN_1938; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1940 = 11'h745 == _T_481 ? _T_6887_1861 : _GEN_1939; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1941 = 11'h746 == _T_481 ? _T_6887_1862 : _GEN_1940; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1942 = 11'h747 == _T_481 ? _T_6887_1863 : _GEN_1941; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1943 = 11'h748 == _T_481 ? _T_6887_1864 : _GEN_1942; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1944 = 11'h749 == _T_481 ? _T_6887_1865 : _GEN_1943; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1945 = 11'h74a == _T_481 ? _T_6887_1866 : _GEN_1944; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1946 = 11'h74b == _T_481 ? _T_6887_1867 : _GEN_1945; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1947 = 11'h74c == _T_481 ? _T_6887_1868 : _GEN_1946; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1948 = 11'h74d == _T_481 ? _T_6887_1869 : _GEN_1947; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1949 = 11'h74e == _T_481 ? _T_6887_1870 : _GEN_1948; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1950 = 11'h74f == _T_481 ? _T_6887_1871 : _GEN_1949; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1951 = 11'h750 == _T_481 ? _T_6887_1872 : _GEN_1950; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1952 = 11'h751 == _T_481 ? _T_6887_1873 : _GEN_1951; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1953 = 11'h752 == _T_481 ? _T_6887_1874 : _GEN_1952; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1954 = 11'h753 == _T_481 ? _T_6887_1875 : _GEN_1953; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1955 = 11'h754 == _T_481 ? _T_6887_1876 : _GEN_1954; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1956 = 11'h755 == _T_481 ? _T_6887_1877 : _GEN_1955; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1957 = 11'h756 == _T_481 ? _T_6887_1878 : _GEN_1956; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1958 = 11'h757 == _T_481 ? _T_6887_1879 : _GEN_1957; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1959 = 11'h758 == _T_481 ? _T_6887_1880 : _GEN_1958; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1960 = 11'h759 == _T_481 ? _T_6887_1881 : _GEN_1959; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1961 = 11'h75a == _T_481 ? _T_6887_1882 : _GEN_1960; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1962 = 11'h75b == _T_481 ? _T_6887_1883 : _GEN_1961; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1963 = 11'h75c == _T_481 ? _T_6887_1884 : _GEN_1962; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1964 = 11'h75d == _T_481 ? _T_6887_1885 : _GEN_1963; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1965 = 11'h75e == _T_481 ? _T_6887_1886 : _GEN_1964; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1966 = 11'h75f == _T_481 ? _T_6887_1887 : _GEN_1965; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1967 = 11'h760 == _T_481 ? _T_6887_1888 : _GEN_1966; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1968 = 11'h761 == _T_481 ? _T_6887_1889 : _GEN_1967; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1969 = 11'h762 == _T_481 ? _T_6887_1890 : _GEN_1968; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1970 = 11'h763 == _T_481 ? _T_6887_1891 : _GEN_1969; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1971 = 11'h764 == _T_481 ? _T_6887_1892 : _GEN_1970; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1972 = 11'h765 == _T_481 ? _T_6887_1893 : _GEN_1971; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1973 = 11'h766 == _T_481 ? _T_6887_1894 : _GEN_1972; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1974 = 11'h767 == _T_481 ? _T_6887_1895 : _GEN_1973; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1975 = 11'h768 == _T_481 ? _T_6887_1896 : _GEN_1974; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1976 = 11'h769 == _T_481 ? _T_6887_1897 : _GEN_1975; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1977 = 11'h76a == _T_481 ? _T_6887_1898 : _GEN_1976; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1978 = 11'h76b == _T_481 ? _T_6887_1899 : _GEN_1977; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1979 = 11'h76c == _T_481 ? _T_6887_1900 : _GEN_1978; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1980 = 11'h76d == _T_481 ? _T_6887_1901 : _GEN_1979; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1981 = 11'h76e == _T_481 ? _T_6887_1902 : _GEN_1980; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1982 = 11'h76f == _T_481 ? _T_6887_1903 : _GEN_1981; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1983 = 11'h770 == _T_481 ? _T_6887_1904 : _GEN_1982; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1984 = 11'h771 == _T_481 ? _T_6887_1905 : _GEN_1983; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1985 = 11'h772 == _T_481 ? _T_6887_1906 : _GEN_1984; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1986 = 11'h773 == _T_481 ? _T_6887_1907 : _GEN_1985; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1987 = 11'h774 == _T_481 ? _T_6887_1908 : _GEN_1986; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1988 = 11'h775 == _T_481 ? _T_6887_1909 : _GEN_1987; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1989 = 11'h776 == _T_481 ? _T_6887_1910 : _GEN_1988; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1990 = 11'h777 == _T_481 ? _T_6887_1911 : _GEN_1989; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1991 = 11'h778 == _T_481 ? _T_6887_1912 : _GEN_1990; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1992 = 11'h779 == _T_481 ? _T_6887_1913 : _GEN_1991; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1993 = 11'h77a == _T_481 ? _T_6887_1914 : _GEN_1992; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1994 = 11'h77b == _T_481 ? _T_6887_1915 : _GEN_1993; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1995 = 11'h77c == _T_481 ? _T_6887_1916 : _GEN_1994; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1996 = 11'h77d == _T_481 ? _T_6887_1917 : _GEN_1995; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1997 = 11'h77e == _T_481 ? _T_6887_1918 : _GEN_1996; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1998 = 11'h77f == _T_481 ? _T_6887_1919 : _GEN_1997; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_1999 = 11'h780 == _T_481 ? _T_6887_1920 : _GEN_1998; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2000 = 11'h781 == _T_481 ? _T_6887_1921 : _GEN_1999; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2001 = 11'h782 == _T_481 ? _T_6887_1922 : _GEN_2000; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2002 = 11'h783 == _T_481 ? _T_6887_1923 : _GEN_2001; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2003 = 11'h784 == _T_481 ? _T_6887_1924 : _GEN_2002; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2004 = 11'h785 == _T_481 ? _T_6887_1925 : _GEN_2003; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2005 = 11'h786 == _T_481 ? _T_6887_1926 : _GEN_2004; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2006 = 11'h787 == _T_481 ? _T_6887_1927 : _GEN_2005; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2007 = 11'h788 == _T_481 ? _T_6887_1928 : _GEN_2006; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2008 = 11'h789 == _T_481 ? _T_6887_1929 : _GEN_2007; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2009 = 11'h78a == _T_481 ? _T_6887_1930 : _GEN_2008; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2010 = 11'h78b == _T_481 ? _T_6887_1931 : _GEN_2009; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2011 = 11'h78c == _T_481 ? _T_6887_1932 : _GEN_2010; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2012 = 11'h78d == _T_481 ? _T_6887_1933 : _GEN_2011; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2013 = 11'h78e == _T_481 ? _T_6887_1934 : _GEN_2012; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2014 = 11'h78f == _T_481 ? _T_6887_1935 : _GEN_2013; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2015 = 11'h790 == _T_481 ? _T_6887_1936 : _GEN_2014; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2016 = 11'h791 == _T_481 ? _T_6887_1937 : _GEN_2015; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2017 = 11'h792 == _T_481 ? _T_6887_1938 : _GEN_2016; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2018 = 11'h793 == _T_481 ? _T_6887_1939 : _GEN_2017; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2019 = 11'h794 == _T_481 ? _T_6887_1940 : _GEN_2018; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2020 = 11'h795 == _T_481 ? _T_6887_1941 : _GEN_2019; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2021 = 11'h796 == _T_481 ? _T_6887_1942 : _GEN_2020; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2022 = 11'h797 == _T_481 ? _T_6887_1943 : _GEN_2021; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2023 = 11'h798 == _T_481 ? _T_6887_1944 : _GEN_2022; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2024 = 11'h799 == _T_481 ? _T_6887_1945 : _GEN_2023; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2025 = 11'h79a == _T_481 ? _T_6887_1946 : _GEN_2024; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2026 = 11'h79b == _T_481 ? _T_6887_1947 : _GEN_2025; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2027 = 11'h79c == _T_481 ? _T_6887_1948 : _GEN_2026; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2028 = 11'h79d == _T_481 ? _T_6887_1949 : _GEN_2027; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2029 = 11'h79e == _T_481 ? _T_6887_1950 : _GEN_2028; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2030 = 11'h79f == _T_481 ? _T_6887_1951 : _GEN_2029; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2031 = 11'h7a0 == _T_481 ? _T_6887_1952 : _GEN_2030; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2032 = 11'h7a1 == _T_481 ? _T_6887_1953 : _GEN_2031; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2033 = 11'h7a2 == _T_481 ? _T_6887_1954 : _GEN_2032; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2034 = 11'h7a3 == _T_481 ? _T_6887_1955 : _GEN_2033; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2035 = 11'h7a4 == _T_481 ? _T_6887_1956 : _GEN_2034; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2036 = 11'h7a5 == _T_481 ? _T_6887_1957 : _GEN_2035; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2037 = 11'h7a6 == _T_481 ? _T_6887_1958 : _GEN_2036; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2038 = 11'h7a7 == _T_481 ? _T_6887_1959 : _GEN_2037; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2039 = 11'h7a8 == _T_481 ? _T_6887_1960 : _GEN_2038; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2040 = 11'h7a9 == _T_481 ? _T_6887_1961 : _GEN_2039; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2041 = 11'h7aa == _T_481 ? _T_6887_1962 : _GEN_2040; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2042 = 11'h7ab == _T_481 ? _T_6887_1963 : _GEN_2041; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2043 = 11'h7ac == _T_481 ? _T_6887_1964 : _GEN_2042; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2044 = 11'h7ad == _T_481 ? _T_6887_1965 : _GEN_2043; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2045 = 11'h7ae == _T_481 ? _T_6887_1966 : _GEN_2044; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2046 = 11'h7af == _T_481 ? _T_6887_1967 : _GEN_2045; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2047 = 11'h7b0 == _T_481 ? _T_6887_1968 : _GEN_2046; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2048 = 11'h7b1 == _T_481 ? _T_6887_1969 : _GEN_2047; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2049 = 11'h7b2 == _T_481 ? _T_6887_1970 : _GEN_2048; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2050 = 11'h7b3 == _T_481 ? _T_6887_1971 : _GEN_2049; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2051 = 11'h7b4 == _T_481 ? _T_6887_1972 : _GEN_2050; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2052 = 11'h7b5 == _T_481 ? _T_6887_1973 : _GEN_2051; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2053 = 11'h7b6 == _T_481 ? _T_6887_1974 : _GEN_2052; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2054 = 11'h7b7 == _T_481 ? _T_6887_1975 : _GEN_2053; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2055 = 11'h7b8 == _T_481 ? _T_6887_1976 : _GEN_2054; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2056 = 11'h7b9 == _T_481 ? _T_6887_1977 : _GEN_2055; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2057 = 11'h7ba == _T_481 ? _T_6887_1978 : _GEN_2056; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2058 = 11'h7bb == _T_481 ? _T_6887_1979 : _GEN_2057; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2059 = 11'h7bc == _T_481 ? _T_6887_1980 : _GEN_2058; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2060 = 11'h7bd == _T_481 ? _T_6887_1981 : _GEN_2059; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2061 = 11'h7be == _T_481 ? _T_6887_1982 : _GEN_2060; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2062 = 11'h7bf == _T_481 ? _T_6887_1983 : _GEN_2061; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2063 = 11'h7c0 == _T_481 ? _T_6887_1984 : _GEN_2062; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2064 = 11'h7c1 == _T_481 ? _T_6887_1985 : _GEN_2063; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2065 = 11'h7c2 == _T_481 ? _T_6887_1986 : _GEN_2064; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2066 = 11'h7c3 == _T_481 ? _T_6887_1987 : _GEN_2065; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2067 = 11'h7c4 == _T_481 ? _T_6887_1988 : _GEN_2066; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2068 = 11'h7c5 == _T_481 ? _T_6887_1989 : _GEN_2067; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2069 = 11'h7c6 == _T_481 ? _T_6887_1990 : _GEN_2068; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2070 = 11'h7c7 == _T_481 ? _T_6887_1991 : _GEN_2069; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2071 = 11'h7c8 == _T_481 ? _T_6887_1992 : _GEN_2070; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2072 = 11'h7c9 == _T_481 ? _T_6887_1993 : _GEN_2071; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2073 = 11'h7ca == _T_481 ? _T_6887_1994 : _GEN_2072; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2074 = 11'h7cb == _T_481 ? _T_6887_1995 : _GEN_2073; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2075 = 11'h7cc == _T_481 ? _T_6887_1996 : _GEN_2074; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2076 = 11'h7cd == _T_481 ? _T_6887_1997 : _GEN_2075; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2077 = 11'h7ce == _T_481 ? _T_6887_1998 : _GEN_2076; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2078 = 11'h7cf == _T_481 ? _T_6887_1999 : _GEN_2077; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2079 = 11'h7d0 == _T_481 ? _T_6887_2000 : _GEN_2078; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2080 = 11'h7d1 == _T_481 ? _T_6887_2001 : _GEN_2079; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2081 = 11'h7d2 == _T_481 ? _T_6887_2002 : _GEN_2080; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2082 = 11'h7d3 == _T_481 ? _T_6887_2003 : _GEN_2081; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2083 = 11'h7d4 == _T_481 ? _T_6887_2004 : _GEN_2082; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2084 = 11'h7d5 == _T_481 ? _T_6887_2005 : _GEN_2083; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2085 = 11'h7d6 == _T_481 ? _T_6887_2006 : _GEN_2084; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2086 = 11'h7d7 == _T_481 ? _T_6887_2007 : _GEN_2085; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2087 = 11'h7d8 == _T_481 ? _T_6887_2008 : _GEN_2086; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2088 = 11'h7d9 == _T_481 ? _T_6887_2009 : _GEN_2087; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2089 = 11'h7da == _T_481 ? _T_6887_2010 : _GEN_2088; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2090 = 11'h7db == _T_481 ? _T_6887_2011 : _GEN_2089; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2091 = 11'h7dc == _T_481 ? _T_6887_2012 : _GEN_2090; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2092 = 11'h7dd == _T_481 ? _T_6887_2013 : _GEN_2091; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2093 = 11'h7de == _T_481 ? _T_6887_2014 : _GEN_2092; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2094 = 11'h7df == _T_481 ? _T_6887_2015 : _GEN_2093; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2095 = 11'h7e0 == _T_481 ? _T_6887_2016 : _GEN_2094; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2096 = 11'h7e1 == _T_481 ? _T_6887_2017 : _GEN_2095; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2097 = 11'h7e2 == _T_481 ? _T_6887_2018 : _GEN_2096; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2098 = 11'h7e3 == _T_481 ? _T_6887_2019 : _GEN_2097; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2099 = 11'h7e4 == _T_481 ? _T_6887_2020 : _GEN_2098; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2100 = 11'h7e5 == _T_481 ? _T_6887_2021 : _GEN_2099; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2101 = 11'h7e6 == _T_481 ? _T_6887_2022 : _GEN_2100; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2102 = 11'h7e7 == _T_481 ? _T_6887_2023 : _GEN_2101; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2103 = 11'h7e8 == _T_481 ? _T_6887_2024 : _GEN_2102; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2104 = 11'h7e9 == _T_481 ? _T_6887_2025 : _GEN_2103; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2105 = 11'h7ea == _T_481 ? _T_6887_2026 : _GEN_2104; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2106 = 11'h7eb == _T_481 ? _T_6887_2027 : _GEN_2105; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2107 = 11'h7ec == _T_481 ? _T_6887_2028 : _GEN_2106; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2108 = 11'h7ed == _T_481 ? _T_6887_2029 : _GEN_2107; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2109 = 11'h7ee == _T_481 ? _T_6887_2030 : _GEN_2108; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2110 = 11'h7ef == _T_481 ? _T_6887_2031 : _GEN_2109; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2111 = 11'h7f0 == _T_481 ? _T_6887_2032 : _GEN_2110; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2112 = 11'h7f1 == _T_481 ? _T_6887_2033 : _GEN_2111; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2113 = 11'h7f2 == _T_481 ? _T_6887_2034 : _GEN_2112; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2114 = 11'h7f3 == _T_481 ? _T_6887_2035 : _GEN_2113; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2115 = 11'h7f4 == _T_481 ? _T_6887_2036 : _GEN_2114; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2116 = 11'h7f5 == _T_481 ? _T_6887_2037 : _GEN_2115; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2117 = 11'h7f6 == _T_481 ? _T_6887_2038 : _GEN_2116; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2118 = 11'h7f7 == _T_481 ? _T_6887_2039 : _GEN_2117; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2119 = 11'h7f8 == _T_481 ? _T_6887_2040 : _GEN_2118; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2120 = 11'h7f9 == _T_481 ? _T_6887_2041 : _GEN_2119; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2121 = 11'h7fa == _T_481 ? _T_6887_2042 : _GEN_2120; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2122 = 11'h7fb == _T_481 ? _T_6887_2043 : _GEN_2121; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2123 = 11'h7fc == _T_481 ? _T_6887_2044 : _GEN_2122; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2124 = 11'h7fd == _T_481 ? _T_6887_2045 : _GEN_2123; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2125 = 11'h7fe == _T_481 ? _T_6887_2046 : _GEN_2124; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_2126 = 11'h7ff == _T_481 ? _T_6887_2047 : _GEN_2125; // @[TLSimpleL2.scala 331:30:freechips.rocketchip.system.DefaultConfig.fir@223417.6]
  assign _GEN_4175 = _T_13036 ? 4'h6 : _GEN_78; // @[TLSimpleL2.scala 326:40:freechips.rocketchip.system.DefaultConfig.fir@223412.4]
  assign _T_604_0 = L2_meta_array_RW0_rdata_0_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221284.4]
  assign _T_604_1 = L2_meta_array_RW0_rdata_1_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221285.4]
  assign _T_604_2 = L2_meta_array_RW0_rdata_2_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221286.4]
  assign _T_604_3 = L2_meta_array_RW0_rdata_3_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221287.4]
  assign _T_604_4 = L2_meta_array_RW0_rdata_4_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221288.4]
  assign _T_604_5 = L2_meta_array_RW0_rdata_5_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221289.4]
  assign _T_604_6 = L2_meta_array_RW0_rdata_6_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221290.4]
  assign _T_604_7 = L2_meta_array_RW0_rdata_7_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221291.4]
  assign _T_604_8 = L2_meta_array_RW0_rdata_8_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221292.4]
  assign _T_604_9 = L2_meta_array_RW0_rdata_9_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221293.4]
  assign _T_604_10 = L2_meta_array_RW0_rdata_10_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221294.4]
  assign _T_604_11 = L2_meta_array_RW0_rdata_11_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221295.4]
  assign _T_604_12 = L2_meta_array_RW0_rdata_12_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221296.4]
  assign _T_604_13 = L2_meta_array_RW0_rdata_13_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221297.4]
  assign _T_604_14 = L2_meta_array_RW0_rdata_14_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221298.4]
  assign _T_604_15 = L2_meta_array_RW0_rdata_15_tag; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221282.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221299.4]
  assign _T_663_0 = L2_meta_array_RW0_rdata_0_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221335.4]
  assign _T_663_1 = L2_meta_array_RW0_rdata_1_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221336.4]
  assign _T_663_2 = L2_meta_array_RW0_rdata_2_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221337.4]
  assign _T_663_3 = L2_meta_array_RW0_rdata_3_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221338.4]
  assign _T_663_4 = L2_meta_array_RW0_rdata_4_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221339.4]
  assign _T_663_5 = L2_meta_array_RW0_rdata_5_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221340.4]
  assign _T_663_6 = L2_meta_array_RW0_rdata_6_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221341.4]
  assign _T_663_7 = L2_meta_array_RW0_rdata_7_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221342.4]
  assign _T_663_8 = L2_meta_array_RW0_rdata_8_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221343.4]
  assign _T_663_9 = L2_meta_array_RW0_rdata_9_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221344.4]
  assign _T_663_10 = L2_meta_array_RW0_rdata_10_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221345.4]
  assign _T_663_11 = L2_meta_array_RW0_rdata_11_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221346.4]
  assign _T_663_12 = L2_meta_array_RW0_rdata_12_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221347.4]
  assign _T_663_13 = L2_meta_array_RW0_rdata_13_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221348.4]
  assign _T_663_14 = L2_meta_array_RW0_rdata_14_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221349.4]
  assign _T_663_15 = L2_meta_array_RW0_rdata_15_dsid; // @[TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221333.4 TLSimpleL2.scala 304:47:freechips.rocketchip.system.DefaultConfig.fir@221350.4]
  assign _T_13044 = _T_291[32:17]; // @[TLSimpleL2.scala 337:21:freechips.rocketchip.system.DefaultConfig.fir@223422.4]
  assign _T_13045 = _T_690_0 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223423.4]
  assign _T_13046 = _T_690_1 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223424.4]
  assign _T_13047 = _T_690_2 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223425.4]
  assign _T_13048 = _T_690_3 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223426.4]
  assign _T_13049 = _T_690_4 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223427.4]
  assign _T_13050 = _T_690_5 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223428.4]
  assign _T_13051 = _T_690_6 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223429.4]
  assign _T_13052 = _T_690_7 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223430.4]
  assign _T_13053 = _T_690_8 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223431.4]
  assign _T_13054 = _T_690_9 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223432.4]
  assign _T_13055 = _T_690_10 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223433.4]
  assign _T_13056 = _T_690_11 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223434.4]
  assign _T_13057 = _T_690_12 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223435.4]
  assign _T_13058 = _T_690_13 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223436.4]
  assign _T_13059 = _T_690_14 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223437.4]
  assign _T_13060 = _T_690_15 == _T_13044; // @[TLSimpleL2.scala 338:60:freechips.rocketchip.system.DefaultConfig.fir@223438.4]
  assign _T_13083 = _T_684[0]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223457.4]
  assign _T_13084 = _T_13045 & _T_13083; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223458.4]
  assign _T_13085 = _T_684[1]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223459.4]
  assign _T_13086 = _T_13046 & _T_13085; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223460.4]
  assign _T_13087 = _T_684[2]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223461.4]
  assign _T_13088 = _T_13047 & _T_13087; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223462.4]
  assign _T_13089 = _T_684[3]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223463.4]
  assign _T_13090 = _T_13048 & _T_13089; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223464.4]
  assign _T_13091 = _T_684[4]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223465.4]
  assign _T_13092 = _T_13049 & _T_13091; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223466.4]
  assign _T_13093 = _T_684[5]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223467.4]
  assign _T_13094 = _T_13050 & _T_13093; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223468.4]
  assign _T_13095 = _T_684[6]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223469.4]
  assign _T_13096 = _T_13051 & _T_13095; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223470.4]
  assign _T_13097 = _T_684[7]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223471.4]
  assign _T_13098 = _T_13052 & _T_13097; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223472.4]
  assign _T_13099 = _T_684[8]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223473.4]
  assign _T_13100 = _T_13053 & _T_13099; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223474.4]
  assign _T_13101 = _T_684[9]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223475.4]
  assign _T_13102 = _T_13054 & _T_13101; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223476.4]
  assign _T_13103 = _T_684[10]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223477.4]
  assign _T_13104 = _T_13055 & _T_13103; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223478.4]
  assign _T_13105 = _T_684[11]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223479.4]
  assign _T_13106 = _T_13056 & _T_13105; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223480.4]
  assign _T_13107 = _T_684[12]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223481.4]
  assign _T_13108 = _T_13057 & _T_13107; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223482.4]
  assign _T_13109 = _T_684[13]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223483.4]
  assign _T_13110 = _T_13058 & _T_13109; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223484.4]
  assign _T_13111 = _T_684[14]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223485.4]
  assign _T_13112 = _T_13059 & _T_13111; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223486.4]
  assign _T_13113 = _T_684[15]; // @[TLSimpleL2.scala 339:75:freechips.rocketchip.system.DefaultConfig.fir@223487.4]
  assign _T_13114 = _T_13060 & _T_13113; // @[TLSimpleL2.scala 339:60:freechips.rocketchip.system.DefaultConfig.fir@223488.4]
  assign _T_13137 = {_T_13086,_T_13084}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223507.4]
  assign _T_13138 = {_T_13090,_T_13088}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223508.4]
  assign _T_13139 = {_T_13138,_T_13137}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223509.4]
  assign _T_13140 = {_T_13094,_T_13092}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223510.4]
  assign _T_13141 = {_T_13098,_T_13096}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223511.4]
  assign _T_13142 = {_T_13141,_T_13140}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223512.4]
  assign _T_13143 = {_T_13142,_T_13139}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223513.4]
  assign _T_13144 = {_T_13102,_T_13100}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223514.4]
  assign _T_13145 = {_T_13106,_T_13104}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223515.4]
  assign _T_13146 = {_T_13145,_T_13144}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223516.4]
  assign _T_13147 = {_T_13110,_T_13108}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223517.4]
  assign _T_13148 = {_T_13114,_T_13112}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223518.4]
  assign _T_13149 = {_T_13148,_T_13147}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223519.4]
  assign _T_13150 = {_T_13149,_T_13146}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223520.4]
  assign _T_13151 = {_T_13150,_T_13143}; // @[TLSimpleL2.scala 339:80:freechips.rocketchip.system.DefaultConfig.fir@223521.4]
  assign _T_13152 = _T_13151 != 16'h0; // @[TLSimpleL2.scala 340:31:freechips.rocketchip.system.DefaultConfig.fir@223522.4]
  assign _T_13153 = _T_13152 & _T_301; // @[TLSimpleL2.scala 341:26:freechips.rocketchip.system.DefaultConfig.fir@223523.4]
  assign _T_13154 = _T_13152 & _T_303; // @[TLSimpleL2.scala 342:27:freechips.rocketchip.system.DefaultConfig.fir@223524.4]
  assign _T_13155 = _T_13152 == 1'h0; // @[TLSimpleL2.scala 343:23:freechips.rocketchip.system.DefaultConfig.fir@223525.4]
  assign _T_13156 = _T_13155 & _T_301; // @[TLSimpleL2.scala 343:28:freechips.rocketchip.system.DefaultConfig.fir@223526.4]
  assign _T_13158 = _T_13155 & _T_303; // @[TLSimpleL2.scala 344:29:freechips.rocketchip.system.DefaultConfig.fir@223528.4]
  assign _T_13162 = _T_13151[1]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223536.4]
  assign _T_13163 = _T_13151[2]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223540.4]
  assign _GEN_6261 = _T_13163 ? 2'h2 : {{1'd0}, _T_13162}; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223541.4]
  assign _T_13164 = _T_13151[3]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223544.4]
  assign _GEN_6262 = _T_13164 ? 2'h3 : _GEN_6261; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223545.4]
  assign _T_13165 = _T_13151[4]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223548.4]
  assign _GEN_6263 = _T_13165 ? 3'h4 : {{1'd0}, _GEN_6262}; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223549.4]
  assign _T_13166 = _T_13151[5]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223552.4]
  assign _GEN_6264 = _T_13166 ? 3'h5 : _GEN_6263; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223553.4]
  assign _T_13167 = _T_13151[6]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223556.4]
  assign _GEN_6265 = _T_13167 ? 3'h6 : _GEN_6264; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223557.4]
  assign _T_13168 = _T_13151[7]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223560.4]
  assign _GEN_6266 = _T_13168 ? 3'h7 : _GEN_6265; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223561.4]
  assign _T_13169 = _T_13151[8]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223564.4]
  assign _GEN_6267 = _T_13169 ? 4'h8 : {{1'd0}, _GEN_6266}; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223565.4]
  assign _T_13170 = _T_13151[9]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223568.4]
  assign _GEN_6268 = _T_13170 ? 4'h9 : _GEN_6267; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223569.4]
  assign _T_13171 = _T_13151[10]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223572.4]
  assign _GEN_6269 = _T_13171 ? 4'ha : _GEN_6268; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223573.4]
  assign _T_13172 = _T_13151[11]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223576.4]
  assign _GEN_6270 = _T_13172 ? 4'hb : _GEN_6269; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223577.4]
  assign _T_13173 = _T_13151[12]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223580.4]
  assign _GEN_6271 = _T_13173 ? 4'hc : _GEN_6270; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223581.4]
  assign _T_13174 = _T_13151[13]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223584.4]
  assign _GEN_6272 = _T_13174 ? 4'hd : _GEN_6271; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223585.4]
  assign _T_13175 = _T_13151[14]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223588.4]
  assign _GEN_6273 = _T_13175 ? 4'he : _GEN_6272; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223589.4]
  assign _T_13176 = _T_13151[15]; // @[TLSimpleL2.scala 347:55:freechips.rocketchip.system.DefaultConfig.fir@223592.4]
  assign _GEN_6274 = _T_13176 ? 4'hf : _GEN_6273; // @[TLSimpleL2.scala 347:60:freechips.rocketchip.system.DefaultConfig.fir@223593.4]
  assign _T_13177 = _T_710 & cp_waymask; // @[TLSimpleL2.scala 351:42:freechips.rocketchip.system.DefaultConfig.fir@223597.4]
  assign _T_13178 = _T_13177 != 16'h0; // @[TLSimpleL2.scala 351:55:freechips.rocketchip.system.DefaultConfig.fir@223598.4]
  assign _T_13180 = _T_13177[0]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223600.4]
  assign _T_13181 = _T_13177[1]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223601.4]
  assign _T_13182 = _T_13177[2]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223602.4]
  assign _T_13183 = _T_13177[3]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223603.4]
  assign _T_13184 = _T_13177[4]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223604.4]
  assign _T_13185 = _T_13177[5]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223605.4]
  assign _T_13186 = _T_13177[6]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223606.4]
  assign _T_13187 = _T_13177[7]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223607.4]
  assign _T_13188 = _T_13177[8]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223608.4]
  assign _T_13189 = _T_13177[9]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223609.4]
  assign _T_13190 = _T_13177[10]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223610.4]
  assign _T_13191 = _T_13177[11]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223611.4]
  assign _T_13192 = _T_13177[12]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223612.4]
  assign _T_13193 = _T_13177[13]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223613.4]
  assign _T_13194 = _T_13177[14]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223614.4]
  assign _T_13196 = _T_13194 ? 4'he : 4'hf; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223616.4]
  assign _T_13197 = _T_13193 ? 4'hd : _T_13196; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223617.4]
  assign _T_13198 = _T_13192 ? 4'hc : _T_13197; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223618.4]
  assign _T_13199 = _T_13191 ? 4'hb : _T_13198; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223619.4]
  assign _T_13200 = _T_13190 ? 4'ha : _T_13199; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223620.4]
  assign _T_13201 = _T_13189 ? 4'h9 : _T_13200; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223621.4]
  assign _T_13202 = _T_13188 ? 4'h8 : _T_13201; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223622.4]
  assign _T_13203 = _T_13187 ? 4'h7 : _T_13202; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223623.4]
  assign _T_13204 = _T_13186 ? 4'h6 : _T_13203; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223624.4]
  assign _T_13205 = _T_13185 ? 4'h5 : _T_13204; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223625.4]
  assign _T_13206 = _T_13184 ? 4'h4 : _T_13205; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223626.4]
  assign _T_13207 = _T_13183 ? 4'h3 : _T_13206; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223627.4]
  assign _T_13208 = _T_13182 ? 4'h2 : _T_13207; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223628.4]
  assign _T_13209 = _T_13181 ? 4'h1 : _T_13208; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223629.4]
  assign _T_13210 = _T_13180 ? 4'h0 : _T_13209; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223630.4]
  assign _T_13211 = cp_waymask != 16'h0; // @[TLSimpleL2.scala 352:23:freechips.rocketchip.system.DefaultConfig.fir@223631.4]
  assign _T_13212 = cp_waymask[0]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223632.4]
  assign _T_13213 = cp_waymask[1]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223633.4]
  assign _T_13214 = cp_waymask[2]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223634.4]
  assign _T_13215 = cp_waymask[3]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223635.4]
  assign _T_13216 = cp_waymask[4]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223636.4]
  assign _T_13217 = cp_waymask[5]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223637.4]
  assign _T_13218 = cp_waymask[6]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223638.4]
  assign _T_13219 = cp_waymask[7]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223639.4]
  assign _T_13220 = cp_waymask[8]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223640.4]
  assign _T_13221 = cp_waymask[9]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223641.4]
  assign _T_13222 = cp_waymask[10]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223642.4]
  assign _T_13223 = cp_waymask[11]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223643.4]
  assign _T_13224 = cp_waymask[12]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223644.4]
  assign _T_13225 = cp_waymask[13]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223645.4]
  assign _T_13226 = cp_waymask[14]; // @[OneHot.scala 39:40:freechips.rocketchip.system.DefaultConfig.fir@223646.4]
  assign _T_13228 = _T_13226 ? 4'he : 4'hf; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223648.4]
  assign _T_13229 = _T_13225 ? 4'hd : _T_13228; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223649.4]
  assign _T_13230 = _T_13224 ? 4'hc : _T_13229; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223650.4]
  assign _T_13231 = _T_13223 ? 4'hb : _T_13230; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223651.4]
  assign _T_13232 = _T_13222 ? 4'ha : _T_13231; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223652.4]
  assign _T_13233 = _T_13221 ? 4'h9 : _T_13232; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223653.4]
  assign _T_13234 = _T_13220 ? 4'h8 : _T_13233; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223654.4]
  assign _T_13235 = _T_13219 ? 4'h7 : _T_13234; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223655.4]
  assign _T_13236 = _T_13218 ? 4'h6 : _T_13235; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223656.4]
  assign _T_13237 = _T_13217 ? 4'h5 : _T_13236; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223657.4]
  assign _T_13238 = _T_13216 ? 4'h4 : _T_13237; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223658.4]
  assign _T_13239 = _T_13215 ? 4'h3 : _T_13238; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223659.4]
  assign _T_13240 = _T_13214 ? 4'h2 : _T_13239; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223660.4]
  assign _T_13241 = _T_13213 ? 4'h1 : _T_13240; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223661.4]
  assign _T_13242 = _T_13212 ? 4'h0 : _T_13241; // @[Mux.scala 31:69:freechips.rocketchip.system.DefaultConfig.fir@223662.4]
  assign _T_13243 = _T_13211 ? _T_13242 : 4'h0; // @[TLSimpleL2.scala 352:12:freechips.rocketchip.system.DefaultConfig.fir@223663.4]
  assign _T_13244 = _T_13178 ? _T_13210 : _T_13243; // @[TLSimpleL2.scala 351:25:freechips.rocketchip.system.DefaultConfig.fir@223664.4]
  assign _GEN_6276 = 4'h1 == cp_capacity_dsid ? _T_13304_1 : _T_13304_0; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6277 = 4'h2 == cp_capacity_dsid ? _T_13304_2 : _GEN_6276; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6278 = 4'h3 == cp_capacity_dsid ? _T_13304_3 : _GEN_6277; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6279 = 4'h4 == cp_capacity_dsid ? _T_13304_4 : _GEN_6278; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6280 = 4'h5 == cp_capacity_dsid ? _T_13304_5 : _GEN_6279; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6281 = 4'h6 == cp_capacity_dsid ? _T_13304_6 : _GEN_6280; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6282 = 4'h7 == cp_capacity_dsid ? _T_13304_7 : _GEN_6281; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6283 = 4'h8 == cp_capacity_dsid ? _T_13304_8 : _GEN_6282; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6284 = 4'h9 == cp_capacity_dsid ? _T_13304_9 : _GEN_6283; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6285 = 4'ha == cp_capacity_dsid ? _T_13304_10 : _GEN_6284; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6286 = 4'hb == cp_capacity_dsid ? _T_13304_11 : _GEN_6285; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6287 = 4'hc == cp_capacity_dsid ? _T_13304_12 : _GEN_6286; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6288 = 4'hd == cp_capacity_dsid ? _T_13304_13 : _GEN_6287; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _GEN_6289 = 4'he == cp_capacity_dsid ? _T_13304_14 : _GEN_6288; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign _T_13367 = _T_684 >> _T_13244; // @[TLSimpleL2.scala 365:40:freechips.rocketchip.system.DefaultConfig.fir@223688.4]
  assign _T_13368 = _T_13367[0]; // @[TLSimpleL2.scala 365:40:freechips.rocketchip.system.DefaultConfig.fir@223689.4]
  assign _T_13369 = _T_686 >> _T_13244; // @[TLSimpleL2.scala 365:66:freechips.rocketchip.system.DefaultConfig.fir@223690.4]
  assign _T_13370 = _T_13369[0]; // @[TLSimpleL2.scala 365:66:freechips.rocketchip.system.DefaultConfig.fir@223691.4]
  assign _T_13371 = _T_13368 & _T_13370; // @[TLSimpleL2.scala 365:51:freechips.rocketchip.system.DefaultConfig.fir@223692.4]
  assign _T_13373 = {_T_481,6'h0}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223693.4]
  assign _GEN_6292 = 4'h1 == _T_13244 ? _T_690_1 : _T_690_0; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6293 = 4'h2 == _T_13244 ? _T_690_2 : _GEN_6292; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6294 = 4'h3 == _T_13244 ? _T_690_3 : _GEN_6293; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6295 = 4'h4 == _T_13244 ? _T_690_4 : _GEN_6294; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6296 = 4'h5 == _T_13244 ? _T_690_5 : _GEN_6295; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6297 = 4'h6 == _T_13244 ? _T_690_6 : _GEN_6296; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6298 = 4'h7 == _T_13244 ? _T_690_7 : _GEN_6297; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6299 = 4'h8 == _T_13244 ? _T_690_8 : _GEN_6298; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6300 = 4'h9 == _T_13244 ? _T_690_9 : _GEN_6299; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6301 = 4'ha == _T_13244 ? _T_690_10 : _GEN_6300; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6302 = 4'hb == _T_13244 ? _T_690_11 : _GEN_6301; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6303 = 4'hc == _T_13244 ? _T_690_12 : _GEN_6302; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6304 = 4'hd == _T_13244 ? _T_690_13 : _GEN_6303; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6305 = 4'he == _T_13244 ? _T_690_14 : _GEN_6304; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _GEN_6306 = 4'hf == _T_13244 ? _T_690_15 : _GEN_6305; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _T_13374 = {_GEN_6306,_T_13373}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@223694.4]
  assign _T_13375 = _T_13156 & _T_13371; // @[TLSimpleL2.scala 369:43:freechips.rocketchip.system.DefaultConfig.fir@223695.4]
  assign _T_13376 = _T_13371 == 1'h0; // @[TLSimpleL2.scala 370:49:freechips.rocketchip.system.DefaultConfig.fir@223696.4]
  assign _T_13377 = _T_13156 & _T_13376; // @[TLSimpleL2.scala 370:46:freechips.rocketchip.system.DefaultConfig.fir@223697.4]
  assign _T_13378 = _T_13158 & _T_13371; // @[TLSimpleL2.scala 371:45:freechips.rocketchip.system.DefaultConfig.fir@223698.4]
  assign _T_13380 = _T_13158 & _T_13376; // @[TLSimpleL2.scala 372:48:freechips.rocketchip.system.DefaultConfig.fir@223700.4]
  assign _T_13381 = _T_13153 | _T_13154; // @[TLSimpleL2.scala 374:37:freechips.rocketchip.system.DefaultConfig.fir@223701.4]
  assign _T_13382 = _T_13381 | _T_13375; // @[TLSimpleL2.scala 374:50:freechips.rocketchip.system.DefaultConfig.fir@223702.4]
  assign _T_13383 = _T_13382 | _T_13378; // @[TLSimpleL2.scala 374:73:freechips.rocketchip.system.DefaultConfig.fir@223703.4]
  assign _T_13385 = _T_310 < 5'h8; // @[TLSimpleL2.scala 395:31:freechips.rocketchip.system.DefaultConfig.fir@223717.6]
  assign _T_13387 = _T_13385 | reset; // @[TLSimpleL2.scala 395:15:freechips.rocketchip.system.DefaultConfig.fir@223719.6]
  assign _T_13388 = _T_13387 == 1'h0; // @[TLSimpleL2.scala 395:15:freechips.rocketchip.system.DefaultConfig.fir@223720.6]
  assign _T_13392 = _T_13377 | _T_13380; // @[TLSimpleL2.scala 399:45:freechips.rocketchip.system.DefaultConfig.fir@223732.8]
  assign _GEN_6307 = _T_13392 ? 4'hd : _GEN_4175; // @[TLSimpleL2.scala 399:73:freechips.rocketchip.system.DefaultConfig.fir@223733.8]
  assign _GEN_6308 = _T_13383 ? 4'h8 : _GEN_6307; // @[TLSimpleL2.scala 397:85:freechips.rocketchip.system.DefaultConfig.fir@223728.6]
  assign _GEN_6309 = _T_482 ? _GEN_6308 : _GEN_4175; // @[TLSimpleL2.scala 376:35:freechips.rocketchip.system.DefaultConfig.fir@223705.4]
  assign _T_13418 = _T_13152 ? _GEN_6274 : _T_13244; // @[TLSimpleL2.scala 419:27:freechips.rocketchip.system.DefaultConfig.fir@223812.4]
  assign _T_13424 = _T_13178 == 1'h0; // @[TLSimpleL2.scala 422:15:freechips.rocketchip.system.DefaultConfig.fir@223819.6]
  assign _T_13425 = _T_710 | cp_waymask; // @[TLSimpleL2.scala 423:40:freechips.rocketchip.system.DefaultConfig.fir@223821.8]
  assign _T_13426 = 16'h1 << _T_13418; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223825.8]
  assign _T_13428 = ~ _T_710; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223827.8]
  assign _T_13429 = _T_13428 | _T_13426; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223828.8]
  assign _T_13430 = ~ _T_13429; // @[TLSimpleL2.scala 425:46:freechips.rocketchip.system.DefaultConfig.fir@223829.8]
  assign _GEN_6310 = _T_13424 ? _T_13425 : _T_13430; // @[TLSimpleL2.scala 422:50:freechips.rocketchip.system.DefaultConfig.fir@223820.6]
  assign _T_13454 = _T_13418 == 4'h0; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223836.4]
  assign _T_13455 = _T_686 >> _T_13418; // @[TLSimpleL2.scala 437:55:freechips.rocketchip.system.DefaultConfig.fir@223839.6]
  assign _T_13456 = _T_13455[0]; // @[TLSimpleL2.scala 437:55:freechips.rocketchip.system.DefaultConfig.fir@223840.6]
  assign _T_13457 = _T_13156 ? 1'h0 : 1'h1; // @[TLSimpleL2.scala 438:16:freechips.rocketchip.system.DefaultConfig.fir@223841.6]
  assign _T_13458 = _T_13153 ? _T_13456 : _T_13457; // @[TLSimpleL2.scala 437:32:freechips.rocketchip.system.DefaultConfig.fir@223842.6]
  assign _T_13460 = _T_686[0]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223850.6]
  assign _GEN_6312 = _T_13454 ? 1'h1 : _T_13083; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  assign _GEN_6313 = _T_13454 ? _T_13458 : _T_13460; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  assign _GEN_6314 = _T_13454 ? _T_13044 : _T_690_0; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  assign _GEN_6315 = _T_13454 ? _T_297 : _T_714_0; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223837.4]
  assign _T_13461 = _GEN_6310[0]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223855.4]
  assign _T_13462 = _T_13418 == 4'h1; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223857.4]
  assign _T_13468 = _T_686[1]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223871.6]
  assign _GEN_6316 = _T_13462 ? 1'h1 : _T_13085; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  assign _GEN_6317 = _T_13462 ? _T_13458 : _T_13468; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  assign _GEN_6318 = _T_13462 ? _T_13044 : _T_690_1; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  assign _GEN_6319 = _T_13462 ? _T_297 : _T_714_1; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223858.4]
  assign _T_13469 = _GEN_6310[1]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223876.4]
  assign _T_13470 = _T_13418 == 4'h2; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223878.4]
  assign _T_13476 = _T_686[2]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223892.6]
  assign _GEN_6320 = _T_13470 ? 1'h1 : _T_13087; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  assign _GEN_6321 = _T_13470 ? _T_13458 : _T_13476; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  assign _GEN_6322 = _T_13470 ? _T_13044 : _T_690_2; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  assign _GEN_6323 = _T_13470 ? _T_297 : _T_714_2; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223879.4]
  assign _T_13477 = _GEN_6310[2]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223897.4]
  assign _T_13478 = _T_13418 == 4'h3; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223899.4]
  assign _T_13484 = _T_686[3]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223913.6]
  assign _GEN_6324 = _T_13478 ? 1'h1 : _T_13089; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  assign _GEN_6325 = _T_13478 ? _T_13458 : _T_13484; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  assign _GEN_6326 = _T_13478 ? _T_13044 : _T_690_3; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  assign _GEN_6327 = _T_13478 ? _T_297 : _T_714_3; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223900.4]
  assign _T_13485 = _GEN_6310[3]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223918.4]
  assign _T_13486 = _T_13418 == 4'h4; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223920.4]
  assign _T_13492 = _T_686[4]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223934.6]
  assign _GEN_6328 = _T_13486 ? 1'h1 : _T_13091; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  assign _GEN_6329 = _T_13486 ? _T_13458 : _T_13492; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  assign _GEN_6330 = _T_13486 ? _T_13044 : _T_690_4; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  assign _GEN_6331 = _T_13486 ? _T_297 : _T_714_4; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223921.4]
  assign _T_13493 = _GEN_6310[4]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223939.4]
  assign _T_13494 = _T_13418 == 4'h5; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223941.4]
  assign _T_13500 = _T_686[5]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223955.6]
  assign _GEN_6332 = _T_13494 ? 1'h1 : _T_13093; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  assign _GEN_6333 = _T_13494 ? _T_13458 : _T_13500; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  assign _GEN_6334 = _T_13494 ? _T_13044 : _T_690_5; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  assign _GEN_6335 = _T_13494 ? _T_297 : _T_714_5; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223942.4]
  assign _T_13501 = _GEN_6310[5]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223960.4]
  assign _T_13502 = _T_13418 == 4'h6; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223962.4]
  assign _T_13508 = _T_686[6]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223976.6]
  assign _GEN_6336 = _T_13502 ? 1'h1 : _T_13095; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  assign _GEN_6337 = _T_13502 ? _T_13458 : _T_13508; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  assign _GEN_6338 = _T_13502 ? _T_13044 : _T_690_6; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  assign _GEN_6339 = _T_13502 ? _T_297 : _T_714_6; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223963.4]
  assign _T_13509 = _GEN_6310[6]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@223981.4]
  assign _T_13510 = _T_13418 == 4'h7; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@223983.4]
  assign _T_13516 = _T_686[7]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@223997.6]
  assign _GEN_6340 = _T_13510 ? 1'h1 : _T_13097; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  assign _GEN_6341 = _T_13510 ? _T_13458 : _T_13516; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  assign _GEN_6342 = _T_13510 ? _T_13044 : _T_690_7; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  assign _GEN_6343 = _T_13510 ? _T_297 : _T_714_7; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@223984.4]
  assign _T_13517 = _GEN_6310[7]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224002.4]
  assign _T_13518 = _T_13418 == 4'h8; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224004.4]
  assign _T_13524 = _T_686[8]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224018.6]
  assign _GEN_6344 = _T_13518 ? 1'h1 : _T_13099; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  assign _GEN_6345 = _T_13518 ? _T_13458 : _T_13524; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  assign _GEN_6346 = _T_13518 ? _T_13044 : _T_690_8; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  assign _GEN_6347 = _T_13518 ? _T_297 : _T_714_8; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224005.4]
  assign _T_13525 = _GEN_6310[8]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224023.4]
  assign _T_13526 = _T_13418 == 4'h9; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224025.4]
  assign _T_13532 = _T_686[9]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224039.6]
  assign _GEN_6348 = _T_13526 ? 1'h1 : _T_13101; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  assign _GEN_6349 = _T_13526 ? _T_13458 : _T_13532; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  assign _GEN_6350 = _T_13526 ? _T_13044 : _T_690_9; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  assign _GEN_6351 = _T_13526 ? _T_297 : _T_714_9; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224026.4]
  assign _T_13533 = _GEN_6310[9]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224044.4]
  assign _T_13534 = _T_13418 == 4'ha; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224046.4]
  assign _T_13540 = _T_686[10]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224060.6]
  assign _GEN_6352 = _T_13534 ? 1'h1 : _T_13103; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  assign _GEN_6353 = _T_13534 ? _T_13458 : _T_13540; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  assign _GEN_6354 = _T_13534 ? _T_13044 : _T_690_10; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  assign _GEN_6355 = _T_13534 ? _T_297 : _T_714_10; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224047.4]
  assign _T_13541 = _GEN_6310[10]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224065.4]
  assign _T_13542 = _T_13418 == 4'hb; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224067.4]
  assign _T_13548 = _T_686[11]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224081.6]
  assign _GEN_6356 = _T_13542 ? 1'h1 : _T_13105; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  assign _GEN_6357 = _T_13542 ? _T_13458 : _T_13548; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  assign _GEN_6358 = _T_13542 ? _T_13044 : _T_690_11; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  assign _GEN_6359 = _T_13542 ? _T_297 : _T_714_11; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224068.4]
  assign _T_13549 = _GEN_6310[11]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224086.4]
  assign _T_13550 = _T_13418 == 4'hc; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224088.4]
  assign _T_13556 = _T_686[12]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224102.6]
  assign _GEN_6360 = _T_13550 ? 1'h1 : _T_13107; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  assign _GEN_6361 = _T_13550 ? _T_13458 : _T_13556; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  assign _GEN_6362 = _T_13550 ? _T_13044 : _T_690_12; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  assign _GEN_6363 = _T_13550 ? _T_297 : _T_714_12; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224089.4]
  assign _T_13557 = _GEN_6310[12]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224107.4]
  assign _T_13558 = _T_13418 == 4'hd; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224109.4]
  assign _T_13564 = _T_686[13]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224123.6]
  assign _GEN_6364 = _T_13558 ? 1'h1 : _T_13109; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  assign _GEN_6365 = _T_13558 ? _T_13458 : _T_13564; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  assign _GEN_6366 = _T_13558 ? _T_13044 : _T_690_13; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  assign _GEN_6367 = _T_13558 ? _T_297 : _T_714_13; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224110.4]
  assign _T_13565 = _GEN_6310[13]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224128.4]
  assign _T_13566 = _T_13418 == 4'he; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224130.4]
  assign _T_13572 = _T_686[14]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224144.6]
  assign _GEN_6368 = _T_13566 ? 1'h1 : _T_13111; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  assign _GEN_6369 = _T_13566 ? _T_13458 : _T_13572; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  assign _GEN_6370 = _T_13566 ? _T_13044 : _T_690_14; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  assign _GEN_6371 = _T_13566 ? _T_297 : _T_714_14; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224131.4]
  assign _T_13573 = _GEN_6310[14]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224149.4]
  assign _T_13574 = _T_13418 == 4'hf; // @[TLSimpleL2.scala 434:40:freechips.rocketchip.system.DefaultConfig.fir@224151.4]
  assign _T_13580 = _T_686[15]; // @[TLSimpleL2.scala 443:41:freechips.rocketchip.system.DefaultConfig.fir@224165.6]
  assign _GEN_6372 = _T_13574 ? 1'h1 : _T_13113; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  assign _GEN_6373 = _T_13574 ? _T_13458 : _T_13580; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  assign _GEN_6374 = _T_13574 ? _T_13044 : _T_690_15; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  assign _GEN_6375 = _T_13574 ? _T_297 : _T_714_15; // @[TLSimpleL2.scala 435:30:freechips.rocketchip.system.DefaultConfig.fir@224152.4]
  assign _T_13581 = _GEN_6310[15]; // @[TLSimpleL2.scala 447:40:freechips.rocketchip.system.DefaultConfig.fir@224170.4]
  assign _T_13583 = _T_262 ? _T_258 : {{2'd0}, _T_481}; // @[TLSimpleL2.scala 455:32:freechips.rocketchip.system.DefaultConfig.fir@224175.4]
  assign _T_13435_0_dsid = {{12'd0}, _GEN_6315}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223845.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223853.6]
  assign _T_13584_0_dsid = _T_262 ? 16'h0 : _T_13435_0_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_1_dsid = {{12'd0}, _GEN_6319}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223866.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223874.6]
  assign _T_13584_1_dsid = _T_262 ? 16'h0 : _T_13435_1_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_2_dsid = {{12'd0}, _GEN_6323}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223887.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223895.6]
  assign _T_13584_2_dsid = _T_262 ? 16'h0 : _T_13435_2_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_3_dsid = {{12'd0}, _GEN_6327}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223908.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223916.6]
  assign _T_13584_3_dsid = _T_262 ? 16'h0 : _T_13435_3_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_4_dsid = {{12'd0}, _GEN_6331}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223929.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223937.6]
  assign _T_13584_4_dsid = _T_262 ? 16'h0 : _T_13435_4_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_5_dsid = {{12'd0}, _GEN_6335}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223950.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223958.6]
  assign _T_13584_5_dsid = _T_262 ? 16'h0 : _T_13435_5_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_6_dsid = {{12'd0}, _GEN_6339}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223971.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@223979.6]
  assign _T_13584_6_dsid = _T_262 ? 16'h0 : _T_13435_6_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_7_dsid = {{12'd0}, _GEN_6343}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@223992.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224000.6]
  assign _T_13584_7_dsid = _T_262 ? 16'h0 : _T_13435_7_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_8_dsid = {{12'd0}, _GEN_6347}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224013.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224021.6]
  assign _T_13584_8_dsid = _T_262 ? 16'h0 : _T_13435_8_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_9_dsid = {{12'd0}, _GEN_6351}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224034.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224042.6]
  assign _T_13584_9_dsid = _T_262 ? 16'h0 : _T_13435_9_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_10_dsid = {{12'd0}, _GEN_6355}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224055.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224063.6]
  assign _T_13584_10_dsid = _T_262 ? 16'h0 : _T_13435_10_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_11_dsid = {{12'd0}, _GEN_6359}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224076.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224084.6]
  assign _T_13584_11_dsid = _T_262 ? 16'h0 : _T_13435_11_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_12_dsid = {{12'd0}, _GEN_6363}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224097.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224105.6]
  assign _T_13584_12_dsid = _T_262 ? 16'h0 : _T_13435_12_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_13_dsid = {{12'd0}, _GEN_6367}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224118.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224126.6]
  assign _T_13584_13_dsid = _T_262 ? 16'h0 : _T_13435_13_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_14_dsid = {{12'd0}, _GEN_6371}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224139.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224147.6]
  assign _T_13584_14_dsid = _T_262 ? 16'h0 : _T_13435_14_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13435_15_dsid = {{12'd0}, _GEN_6375}; // @[TLSimpleL2.scala 431:33:freechips.rocketchip.system.DefaultConfig.fir@223834.4 TLSimpleL2.scala 440:25:freechips.rocketchip.system.DefaultConfig.fir@224160.6 TLSimpleL2.scala 445:25:freechips.rocketchip.system.DefaultConfig.fir@224168.6]
  assign _T_13584_15_dsid = _T_262 ? 16'h0 : _T_13435_15_dsid; // @[TLSimpleL2.scala 456:33:freechips.rocketchip.system.DefaultConfig.fir@224176.4]
  assign _T_13620 = _T_13583[10:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224178.6]
  assign _T_13659 = _T_13155 & _T_336; // @[TLSimpleL2.scala 461:20:freechips.rocketchip.system.DefaultConfig.fir@224183.6]
  assign _T_13660 = _T_13418 == _T_13244; // @[TLSimpleL2.scala 462:29:freechips.rocketchip.system.DefaultConfig.fir@224185.8]
  assign _T_13662 = _T_13660 | reset; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224187.8]
  assign _T_13663 = _T_13662 == 1'h0; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224188.8]
  assign _T_13666 = 4'h0 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224195.8]
  assign _T_13667 = _T_13368 == 1'h0; // @[TLSimpleL2.scala 465:38:freechips.rocketchip.system.DefaultConfig.fir@224196.8]
  assign _GEN_6377 = 4'h1 == _T_13244 ? _T_714_1 : _T_714_0; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6378 = 4'h2 == _T_13244 ? _T_714_2 : _GEN_6377; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6379 = 4'h3 == _T_13244 ? _T_714_3 : _GEN_6378; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6380 = 4'h4 == _T_13244 ? _T_714_4 : _GEN_6379; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6381 = 4'h5 == _T_13244 ? _T_714_5 : _GEN_6380; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6382 = 4'h6 == _T_13244 ? _T_714_6 : _GEN_6381; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6383 = 4'h7 == _T_13244 ? _T_714_7 : _GEN_6382; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6384 = 4'h8 == _T_13244 ? _T_714_8 : _GEN_6383; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6385 = 4'h9 == _T_13244 ? _T_714_9 : _GEN_6384; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6386 = 4'ha == _T_13244 ? _T_714_10 : _GEN_6385; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6387 = 4'hb == _T_13244 ? _T_714_11 : _GEN_6386; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6388 = 4'hc == _T_13244 ? _T_714_12 : _GEN_6387; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6389 = 4'hd == _T_13244 ? _T_714_13 : _GEN_6388; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6390 = 4'he == _T_13244 ? _T_714_14 : _GEN_6389; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _GEN_6391 = 4'hf == _T_13244 ? _T_714_15 : _GEN_6390; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _T_13668 = 4'h0 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224197.8]
  assign _T_13669 = _T_13667 | _T_13668; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224198.8]
  assign _T_13670 = _T_13666 & _T_13669; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224199.8]
  assign _GEN_6393 = 4'h1 == _T_297 ? _T_13304_1 : _T_13304_0; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6394 = 4'h2 == _T_297 ? _T_13304_2 : _GEN_6393; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6395 = 4'h3 == _T_297 ? _T_13304_3 : _GEN_6394; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6396 = 4'h4 == _T_297 ? _T_13304_4 : _GEN_6395; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6397 = 4'h5 == _T_297 ? _T_13304_5 : _GEN_6396; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6398 = 4'h6 == _T_297 ? _T_13304_6 : _GEN_6397; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6399 = 4'h7 == _T_297 ? _T_13304_7 : _GEN_6398; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6400 = 4'h8 == _T_297 ? _T_13304_8 : _GEN_6399; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6401 = 4'h9 == _T_297 ? _T_13304_9 : _GEN_6400; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6402 = 4'ha == _T_297 ? _T_13304_10 : _GEN_6401; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6403 = 4'hb == _T_297 ? _T_13304_11 : _GEN_6402; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6404 = 4'hc == _T_297 ? _T_13304_12 : _GEN_6403; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6405 = 4'hd == _T_297 ? _T_13304_13 : _GEN_6404; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6406 = 4'he == _T_297 ? _T_13304_14 : _GEN_6405; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _GEN_6407 = 4'hf == _T_297 ? _T_13304_15 : _GEN_6406; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224201.10]
  assign _T_13672 = _GEN_6407 + 15'h1; // @[TLSimpleL2.scala 466:48:freechips.rocketchip.system.DefaultConfig.fir@224202.10]
  assign _T_13673 = 4'h0 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224206.10]
  assign _T_13674 = 4'h0 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224207.10]
  assign _T_13675 = _T_13673 & _T_13674; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224208.10]
  assign _T_13676 = _T_13675 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224209.10]
  assign _GEN_6409 = 4'h1 == _GEN_6391 ? _T_13304_1 : _T_13304_0; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6410 = 4'h2 == _GEN_6391 ? _T_13304_2 : _GEN_6409; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6411 = 4'h3 == _GEN_6391 ? _T_13304_3 : _GEN_6410; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6412 = 4'h4 == _GEN_6391 ? _T_13304_4 : _GEN_6411; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6413 = 4'h5 == _GEN_6391 ? _T_13304_5 : _GEN_6412; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6414 = 4'h6 == _GEN_6391 ? _T_13304_6 : _GEN_6413; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6415 = 4'h7 == _GEN_6391 ? _T_13304_7 : _GEN_6414; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6416 = 4'h8 == _GEN_6391 ? _T_13304_8 : _GEN_6415; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6417 = 4'h9 == _GEN_6391 ? _T_13304_9 : _GEN_6416; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6418 = 4'ha == _GEN_6391 ? _T_13304_10 : _GEN_6417; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6419 = 4'hb == _GEN_6391 ? _T_13304_11 : _GEN_6418; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6420 = 4'hc == _GEN_6391 ? _T_13304_12 : _GEN_6419; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6421 = 4'hd == _GEN_6391 ? _T_13304_13 : _GEN_6420; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6422 = 4'he == _GEN_6391 ? _T_13304_14 : _GEN_6421; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _GEN_6423 = 4'hf == _GEN_6391 ? _T_13304_15 : _GEN_6422; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _T_13677 = _GEN_6423 - 15'h1; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224211.12]
  assign _T_13678 = $unsigned(_T_13677); // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224212.12]
  assign _T_13679 = _T_13678[14:0]; // @[TLSimpleL2.scala 468:45:freechips.rocketchip.system.DefaultConfig.fir@224213.12]
  assign _T_13680 = 4'h1 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224216.8]
  assign _T_13682 = 4'h1 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224218.8]
  assign _T_13683 = _T_13667 | _T_13682; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224219.8]
  assign _T_13684 = _T_13680 & _T_13683; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224220.8]
  assign _T_13687 = 4'h1 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224227.10]
  assign _T_13688 = 4'h1 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224228.10]
  assign _T_13689 = _T_13687 & _T_13688; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224229.10]
  assign _T_13690 = _T_13689 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224230.10]
  assign _T_13694 = 4'h2 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224237.8]
  assign _T_13696 = 4'h2 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224239.8]
  assign _T_13697 = _T_13667 | _T_13696; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224240.8]
  assign _T_13698 = _T_13694 & _T_13697; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224241.8]
  assign _T_13701 = 4'h2 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224248.10]
  assign _T_13702 = 4'h2 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224249.10]
  assign _T_13703 = _T_13701 & _T_13702; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224250.10]
  assign _T_13704 = _T_13703 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224251.10]
  assign _T_13708 = 4'h3 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224258.8]
  assign _T_13710 = 4'h3 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224260.8]
  assign _T_13711 = _T_13667 | _T_13710; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224261.8]
  assign _T_13712 = _T_13708 & _T_13711; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224262.8]
  assign _T_13715 = 4'h3 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224269.10]
  assign _T_13716 = 4'h3 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224270.10]
  assign _T_13717 = _T_13715 & _T_13716; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224271.10]
  assign _T_13718 = _T_13717 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224272.10]
  assign _T_13722 = 4'h4 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224279.8]
  assign _T_13724 = 4'h4 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224281.8]
  assign _T_13725 = _T_13667 | _T_13724; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224282.8]
  assign _T_13726 = _T_13722 & _T_13725; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224283.8]
  assign _T_13729 = 4'h4 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224290.10]
  assign _T_13730 = 4'h4 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224291.10]
  assign _T_13731 = _T_13729 & _T_13730; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224292.10]
  assign _T_13732 = _T_13731 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224293.10]
  assign _T_13736 = 4'h5 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224300.8]
  assign _T_13738 = 4'h5 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224302.8]
  assign _T_13739 = _T_13667 | _T_13738; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224303.8]
  assign _T_13740 = _T_13736 & _T_13739; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224304.8]
  assign _T_13743 = 4'h5 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224311.10]
  assign _T_13744 = 4'h5 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224312.10]
  assign _T_13745 = _T_13743 & _T_13744; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224313.10]
  assign _T_13746 = _T_13745 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224314.10]
  assign _T_13750 = 4'h6 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224321.8]
  assign _T_13752 = 4'h6 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224323.8]
  assign _T_13753 = _T_13667 | _T_13752; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224324.8]
  assign _T_13754 = _T_13750 & _T_13753; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224325.8]
  assign _T_13757 = 4'h6 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224332.10]
  assign _T_13758 = 4'h6 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224333.10]
  assign _T_13759 = _T_13757 & _T_13758; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224334.10]
  assign _T_13760 = _T_13759 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224335.10]
  assign _T_13764 = 4'h7 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224342.8]
  assign _T_13766 = 4'h7 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224344.8]
  assign _T_13767 = _T_13667 | _T_13766; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224345.8]
  assign _T_13768 = _T_13764 & _T_13767; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224346.8]
  assign _T_13771 = 4'h7 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224353.10]
  assign _T_13772 = 4'h7 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224354.10]
  assign _T_13773 = _T_13771 & _T_13772; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224355.10]
  assign _T_13774 = _T_13773 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224356.10]
  assign _T_13778 = 4'h8 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224363.8]
  assign _T_13780 = 4'h8 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224365.8]
  assign _T_13781 = _T_13667 | _T_13780; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224366.8]
  assign _T_13782 = _T_13778 & _T_13781; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224367.8]
  assign _T_13785 = 4'h8 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224374.10]
  assign _T_13786 = 4'h8 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224375.10]
  assign _T_13787 = _T_13785 & _T_13786; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224376.10]
  assign _T_13788 = _T_13787 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224377.10]
  assign _T_13792 = 4'h9 == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224384.8]
  assign _T_13794 = 4'h9 != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224386.8]
  assign _T_13795 = _T_13667 | _T_13794; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224387.8]
  assign _T_13796 = _T_13792 & _T_13795; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224388.8]
  assign _T_13799 = 4'h9 != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224395.10]
  assign _T_13800 = 4'h9 == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224396.10]
  assign _T_13801 = _T_13799 & _T_13800; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224397.10]
  assign _T_13802 = _T_13801 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224398.10]
  assign _T_13806 = 4'ha == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224405.8]
  assign _T_13808 = 4'ha != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224407.8]
  assign _T_13809 = _T_13667 | _T_13808; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224408.8]
  assign _T_13810 = _T_13806 & _T_13809; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224409.8]
  assign _T_13813 = 4'ha != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224416.10]
  assign _T_13814 = 4'ha == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224417.10]
  assign _T_13815 = _T_13813 & _T_13814; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224418.10]
  assign _T_13816 = _T_13815 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224419.10]
  assign _T_13820 = 4'hb == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224426.8]
  assign _T_13822 = 4'hb != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224428.8]
  assign _T_13823 = _T_13667 | _T_13822; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224429.8]
  assign _T_13824 = _T_13820 & _T_13823; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224430.8]
  assign _T_13827 = 4'hb != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224437.10]
  assign _T_13828 = 4'hb == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224438.10]
  assign _T_13829 = _T_13827 & _T_13828; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224439.10]
  assign _T_13830 = _T_13829 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224440.10]
  assign _T_13834 = 4'hc == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224447.8]
  assign _T_13836 = 4'hc != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224449.8]
  assign _T_13837 = _T_13667 | _T_13836; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224450.8]
  assign _T_13838 = _T_13834 & _T_13837; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224451.8]
  assign _T_13841 = 4'hc != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224458.10]
  assign _T_13842 = 4'hc == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224459.10]
  assign _T_13843 = _T_13841 & _T_13842; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224460.10]
  assign _T_13844 = _T_13843 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224461.10]
  assign _T_13848 = 4'hd == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224468.8]
  assign _T_13850 = 4'hd != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224470.8]
  assign _T_13851 = _T_13667 | _T_13850; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224471.8]
  assign _T_13852 = _T_13848 & _T_13851; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224472.8]
  assign _T_13855 = 4'hd != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224479.10]
  assign _T_13856 = 4'hd == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224480.10]
  assign _T_13857 = _T_13855 & _T_13856; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224481.10]
  assign _T_13858 = _T_13857 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224482.10]
  assign _T_13862 = 4'he == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224489.8]
  assign _T_13864 = 4'he != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224491.8]
  assign _T_13865 = _T_13667 | _T_13864; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224492.8]
  assign _T_13866 = _T_13862 & _T_13865; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224493.8]
  assign _T_13869 = 4'he != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224500.10]
  assign _T_13870 = 4'he == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224501.10]
  assign _T_13871 = _T_13869 & _T_13870; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224502.10]
  assign _T_13872 = _T_13871 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224503.10]
  assign _T_13876 = 4'hf == _T_297; // @[TLSimpleL2.scala 465:25:freechips.rocketchip.system.DefaultConfig.fir@224510.8]
  assign _T_13878 = 4'hf != _GEN_6391; // @[TLSimpleL2.scala 465:59:freechips.rocketchip.system.DefaultConfig.fir@224512.8]
  assign _T_13879 = _T_13667 | _T_13878; // @[TLSimpleL2.scala 465:52:freechips.rocketchip.system.DefaultConfig.fir@224513.8]
  assign _T_13880 = _T_13876 & _T_13879; // @[TLSimpleL2.scala 465:34:freechips.rocketchip.system.DefaultConfig.fir@224514.8]
  assign _T_13883 = 4'hf != _T_297; // @[TLSimpleL2.scala 467:30:freechips.rocketchip.system.DefaultConfig.fir@224521.10]
  assign _T_13884 = 4'hf == _GEN_6391; // @[TLSimpleL2.scala 467:46:freechips.rocketchip.system.DefaultConfig.fir@224522.10]
  assign _T_13885 = _T_13883 & _T_13884; // @[TLSimpleL2.scala 467:39:freechips.rocketchip.system.DefaultConfig.fir@224523.10]
  assign _T_13886 = _T_13885 & _T_13368; // @[TLSimpleL2.scala 467:60:freechips.rocketchip.system.DefaultConfig.fir@224524.10]
  assign _T_13891 = _T_13381 ? _GEN_6274 : _T_13244; // @[TLSimpleL2.scala 481:30:freechips.rocketchip.system.DefaultConfig.fir@224536.4]
  assign _T_13895 = _T_482 & _T_13383; // @[TLSimpleL2.scala 484:51:freechips.rocketchip.system.DefaultConfig.fir@224539.4]
  assign _T_13896 = _T_267 == 4'h8; // @[TLSimpleL2.scala 484:80:freechips.rocketchip.system.DefaultConfig.fir@224540.4]
  assign _T_13897 = _T_13893 != 4'h8; // @[TLSimpleL2.scala 484:113:freechips.rocketchip.system.DefaultConfig.fir@224541.4]
  assign _T_13898 = _T_13896 & _T_13897; // @[TLSimpleL2.scala 484:96:freechips.rocketchip.system.DefaultConfig.fir@224542.4]
  assign _T_13899 = _T_13895 | _T_13898; // @[TLSimpleL2.scala 484:70:freechips.rocketchip.system.DefaultConfig.fir@224543.4]
  assign _GEN_7028 = {{3'd0}, _T_481}; // @[TLSimpleL2.scala 485:31:freechips.rocketchip.system.DefaultConfig.fir@224544.4]
  assign _T_13900 = _GEN_7028 << 3; // @[TLSimpleL2.scala 485:31:freechips.rocketchip.system.DefaultConfig.fir@224544.4]
  assign _GEN_7029 = {{10'd0}, _T_13893}; // @[TLSimpleL2.scala 485:59:freechips.rocketchip.system.DefaultConfig.fir@224545.4]
  assign _T_13901 = _T_13900 | _GEN_7029; // @[TLSimpleL2.scala 485:59:freechips.rocketchip.system.DefaultConfig.fir@224545.4]
  assign _T_13909 = _T_13154 ? _GEN_6274 : _T_13244; // @[TLSimpleL2.scala 488:31:freechips.rocketchip.system.DefaultConfig.fir@224548.4]
  assign _T_13912 = _T_267 == 4'h9; // @[TLSimpleL2.scala 490:36:freechips.rocketchip.system.DefaultConfig.fir@224551.4]
  assign _GEN_7031 = {{11'd0}, value_1}; // @[TLSimpleL2.scala 491:60:freechips.rocketchip.system.DefaultConfig.fir@224553.4]
  assign _T_13914 = _T_13900 | _GEN_7031; // @[TLSimpleL2.scala 491:60:freechips.rocketchip.system.DefaultConfig.fir@224553.4]
  assign _T_14156 = {{1'd0}, value_1}; // @[TLSimpleL2.scala 559:49:freechips.rocketchip.system.DefaultConfig.fir@224767.4]
  assign _T_14157 = _T_14156[2:0]; // @[TLSimpleL2.scala 559:49:freechips.rocketchip.system.DefaultConfig.fir@224768.4]
  assign _GEN_6968 = 3'h1 == _T_14157 ? _T_14075_1 : _T_14075_0; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  assign _GEN_6969 = 3'h2 == _T_14157 ? _T_14075_2 : _GEN_6968; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  assign _GEN_6970 = 3'h3 == _T_14157 ? _T_14075_3 : _GEN_6969; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  assign _GEN_6971 = 3'h4 == _T_14157 ? _T_14075_4 : _GEN_6970; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  assign _GEN_6972 = 3'h5 == _T_14157 ? _T_14075_5 : _GEN_6971; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  assign _GEN_6973 = 3'h6 == _T_14157 ? _T_14075_6 : _GEN_6972; // @[TLSimpleL2.scala 560:16:freechips.rocketchip.system.DefaultConfig.fir@224771.4]
  assign _T_14020 = _T_13912 == 1'h0; // @[TLSimpleL2.scala 506:70:freechips.rocketchip.system.DefaultConfig.fir@224644.4]
  assign _T_14021 = _T_13899 & _T_14020; // @[TLSimpleL2.scala 506:67:freechips.rocketchip.system.DefaultConfig.fir@224645.4]
  assign _GEN_6883 = L2_data_array_RW0_rdata_0; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6884 = 4'h1 == _T_13891 ? L2_data_array_RW0_rdata_1 : _GEN_6883; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6885 = 4'h2 == _T_13891 ? L2_data_array_RW0_rdata_2 : _GEN_6884; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6886 = 4'h3 == _T_13891 ? L2_data_array_RW0_rdata_3 : _GEN_6885; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6887 = 4'h4 == _T_13891 ? L2_data_array_RW0_rdata_4 : _GEN_6886; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6888 = 4'h5 == _T_13891 ? L2_data_array_RW0_rdata_5 : _GEN_6887; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6889 = 4'h6 == _T_13891 ? L2_data_array_RW0_rdata_6 : _GEN_6888; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6890 = 4'h7 == _T_13891 ? L2_data_array_RW0_rdata_7 : _GEN_6889; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6891 = 4'h8 == _T_13891 ? L2_data_array_RW0_rdata_8 : _GEN_6890; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6892 = 4'h9 == _T_13891 ? L2_data_array_RW0_rdata_9 : _GEN_6891; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6893 = 4'ha == _T_13891 ? L2_data_array_RW0_rdata_10 : _GEN_6892; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6894 = 4'hb == _T_13891 ? L2_data_array_RW0_rdata_11 : _GEN_6893; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6895 = 4'hc == _T_13891 ? L2_data_array_RW0_rdata_12 : _GEN_6894; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6896 = 4'hd == _T_13891 ? L2_data_array_RW0_rdata_13 : _GEN_6895; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6897 = 4'he == _T_13891 ? L2_data_array_RW0_rdata_14 : _GEN_6896; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _GEN_6898 = 4'hf == _T_13891 ? L2_data_array_RW0_rdata_15 : _GEN_6897; // @[TLSimpleL2.scala 506:17:freechips.rocketchip.system.DefaultConfig.fir@224657.4]
  assign _T_14087 = _T_13893 + 4'h1; // @[TLSimpleL2.scala 517:40:freechips.rocketchip.system.DefaultConfig.fir@224669.6]
  assign _T_14089 = _T_13893 - 4'h1; // @[TLSimpleL2.scala 521:36:freechips.rocketchip.system.DefaultConfig.fir@224674.6]
  assign _T_14090 = $unsigned(_T_14089); // @[TLSimpleL2.scala 521:36:freechips.rocketchip.system.DefaultConfig.fir@224675.6]
  assign _T_14091 = _T_14090[3:0]; // @[TLSimpleL2.scala 521:36:freechips.rocketchip.system.DefaultConfig.fir@224676.6]
  assign _T_14093 = {{1'd0}, _T_14091}; // @[TLSimpleL2.scala 521:57:freechips.rocketchip.system.DefaultConfig.fir@224678.6]
  assign _T_14094 = _T_14093[3:0]; // @[TLSimpleL2.scala 521:57:freechips.rocketchip.system.DefaultConfig.fir@224679.6]
  assign _T_14096 = _T_14094[2:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224680.6]
  assign _T_14097 = _T_13893 == 4'h8; // @[TLSimpleL2.scala 523:29:freechips.rocketchip.system.DefaultConfig.fir@224682.6]
  assign _T_14098 = _T_13375 | _T_13378; // @[TLSimpleL2.scala 527:44:freechips.rocketchip.system.DefaultConfig.fir@224689.10]
  assign _GEN_6908 = _T_13154 ? 4'h7 : _GEN_6309; // @[TLSimpleL2.scala 529:35:freechips.rocketchip.system.DefaultConfig.fir@224694.12]
  assign _GEN_6909 = _T_14098 ? 4'ha : _GEN_6908; // @[TLSimpleL2.scala 527:69:freechips.rocketchip.system.DefaultConfig.fir@224690.10]
  assign _GEN_6910 = _T_13153 ? 4'hf : _GEN_6909; // @[TLSimpleL2.scala 525:27:freechips.rocketchip.system.DefaultConfig.fir@224685.8]
  assign _GEN_6912 = _T_14097 ? _GEN_6910 : _GEN_6309; // @[TLSimpleL2.scala 523:51:freechips.rocketchip.system.DefaultConfig.fir@224683.6]
  assign _GEN_6922 = _T_13896 ? _GEN_6912 : _GEN_6309; // @[TLSimpleL2.scala 519:36:freechips.rocketchip.system.DefaultConfig.fir@224673.4]
  assign _T_14102 = _T_267 == 4'h7; // @[TLSimpleL2.scala 544:19:freechips.rocketchip.system.DefaultConfig.fir@224708.4]
  assign _T_14104 = _T_317 + 3'h1; // @[TLSimpleL2.scala 545:44:freechips.rocketchip.system.DefaultConfig.fir@224711.6]
  assign _T_14106 = {{1'd0}, _T_317}; // @[TLSimpleL2.scala 547:52:freechips.rocketchip.system.DefaultConfig.fir@224714.6]
  assign _T_14107 = _T_14106[2:0]; // @[TLSimpleL2.scala 547:52:freechips.rocketchip.system.DefaultConfig.fir@224715.6]
  assign _GEN_6924 = 3'h1 == _T_14107 ? _T_397_1 : _T_397_0; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _GEN_6925 = 3'h2 == _T_14107 ? _T_397_2 : _GEN_6924; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _GEN_6926 = 3'h3 == _T_14107 ? _T_397_3 : _GEN_6925; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _GEN_6927 = 3'h4 == _T_14107 ? _T_397_4 : _GEN_6926; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _GEN_6928 = 3'h5 == _T_14107 ? _T_397_5 : _GEN_6927; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _GEN_6929 = 3'h6 == _T_14107 ? _T_397_6 : _GEN_6928; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _GEN_6930 = 3'h7 == _T_14107 ? _T_397_7 : _GEN_6929; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _T_14114 = _GEN_6930[0]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224716.6]
  assign _T_14115 = _GEN_6930[1]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224717.6]
  assign _T_14116 = _GEN_6930[2]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224718.6]
  assign _T_14117 = _GEN_6930[3]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224719.6]
  assign _T_14118 = _GEN_6930[4]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224720.6]
  assign _T_14119 = _GEN_6930[5]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224721.6]
  assign _T_14120 = _GEN_6930[6]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224722.6]
  assign _T_14121 = _GEN_6930[7]; // @[Bitwise.scala 27:51:freechips.rocketchip.system.DefaultConfig.fir@224723.6]
  assign _T_14123 = _T_14114 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224725.6]
  assign _T_14125 = _T_14115 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224727.6]
  assign _T_14127 = _T_14116 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224729.6]
  assign _T_14129 = _T_14117 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224731.6]
  assign _T_14131 = _T_14118 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224733.6]
  assign _T_14133 = _T_14119 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224735.6]
  assign _T_14135 = _T_14120 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224737.6]
  assign _T_14137 = _T_14121 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12:freechips.rocketchip.system.DefaultConfig.fir@224739.6]
  assign _T_14138 = {_T_14125,_T_14123}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224740.6]
  assign _T_14139 = {_T_14129,_T_14127}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224741.6]
  assign _T_14140 = {_T_14139,_T_14138}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224742.6]
  assign _T_14141 = {_T_14133,_T_14131}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224743.6]
  assign _T_14142 = {_T_14137,_T_14135}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224744.6]
  assign _T_14143 = {_T_14142,_T_14141}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224745.6]
  assign _T_14144 = {_T_14143,_T_14140}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224746.6]
  assign _T_14145 = ~ _T_14144; // @[TLSimpleL2.scala 542:13:freechips.rocketchip.system.DefaultConfig.fir@224747.6]
  assign _GEN_6932 = 3'h1 == _T_14107 ? _T_14075_1 : _T_14075_0; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6933 = 3'h2 == _T_14107 ? _T_14075_2 : _GEN_6932; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6934 = 3'h3 == _T_14107 ? _T_14075_3 : _GEN_6933; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6935 = 3'h4 == _T_14107 ? _T_14075_4 : _GEN_6934; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6936 = 3'h5 == _T_14107 ? _T_14075_5 : _GEN_6935; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6937 = 3'h6 == _T_14107 ? _T_14075_6 : _GEN_6936; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6938 = 3'h7 == _T_14107 ? _T_14075_7 : _GEN_6937; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _T_14146 = _T_14145 & _GEN_6938; // @[TLSimpleL2.scala 542:25:freechips.rocketchip.system.DefaultConfig.fir@224748.6]
  assign _GEN_6940 = 3'h1 == _T_14107 ? _T_344_1 : _T_344_0; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _GEN_6941 = 3'h2 == _T_14107 ? _T_344_2 : _GEN_6940; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _GEN_6942 = 3'h3 == _T_14107 ? _T_344_3 : _GEN_6941; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _GEN_6943 = 3'h4 == _T_14107 ? _T_344_4 : _GEN_6942; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _GEN_6944 = 3'h5 == _T_14107 ? _T_344_5 : _GEN_6943; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _GEN_6945 = 3'h6 == _T_14107 ? _T_344_6 : _GEN_6944; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _GEN_6946 = 3'h7 == _T_14107 ? _T_344_7 : _GEN_6945; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _T_14147 = _T_14144 & _GEN_6946; // @[TLSimpleL2.scala 542:51:freechips.rocketchip.system.DefaultConfig.fir@224749.6]
  assign _T_14148 = _T_14146 | _T_14147; // @[TLSimpleL2.scala 542:37:freechips.rocketchip.system.DefaultConfig.fir@224750.6]
  assign _GEN_6955 = _T_318 ? 4'h9 : _GEN_6922; // @[TLSimpleL2.scala 550:32:freechips.rocketchip.system.DefaultConfig.fir@224752.6]
  assign _GEN_6965 = _T_14102 ? _GEN_6955 : _GEN_6922; // @[TLSimpleL2.scala 544:41:freechips.rocketchip.system.DefaultConfig.fir@224709.4]
  assign _T_14151 = value_1 == 3'h7; // @[Counter.scala 34:24:freechips.rocketchip.system.DefaultConfig.fir@224759.6]
  assign _T_14153 = value_1 + 3'h1; // @[Counter.scala 35:22:freechips.rocketchip.system.DefaultConfig.fir@224761.6]
  assign _T_14154 = _T_13912 & _T_14151; // @[Counter.scala 64:20:freechips.rocketchip.system.DefaultConfig.fir@224764.4]
  assign _T_14162 = _T_13912 & _T_14154; // @[TLSimpleL2.scala 562:36:freechips.rocketchip.system.DefaultConfig.fir@224773.4]
  assign _GEN_6975 = _T_301 ? 4'hf : 4'h0; // @[TLSimpleL2.scala 563:20:freechips.rocketchip.system.DefaultConfig.fir@224775.6]
  assign _GEN_6976 = _T_14162 ? _GEN_6975 : _GEN_6965; // @[TLSimpleL2.scala 562:51:freechips.rocketchip.system.DefaultConfig.fir@224774.4]
  assign _T_14163 = _T_291[32:6]; // @[TLSimpleL2.scala 574:30:freechips.rocketchip.system.DefaultConfig.fir@224782.4]
  assign _T_14164 = {_T_14163,6'h0}; // @[Cat.scala 30:58:freechips.rocketchip.system.DefaultConfig.fir@224783.4]
  assign _T_14268 = _T_267 == 4'he; // @[TLSimpleL2.scala 647:29:freechips.rocketchip.system.DefaultConfig.fir@224932.4]
  assign _T_14269 = _T_267 == 4'hc; // @[TLSimpleL2.scala 647:58:freechips.rocketchip.system.DefaultConfig.fir@224933.4]
  assign _T_14270 = _T_14268 | _T_14269; // @[TLSimpleL2.scala 647:48:freechips.rocketchip.system.DefaultConfig.fir@224934.4]
  assign _T_14168 = _T_14270 & auto_out_d_valid; // @[Decoupled.scala 37:37:freechips.rocketchip.system.DefaultConfig.fir@224787.4]
  assign _T_14170 = _T_267 == 4'ha; // @[TLSimpleL2.scala 586:19:freechips.rocketchip.system.DefaultConfig.fir@224789.4]
  assign _GEN_6977 = _T_14170 ? 4'hb : _GEN_6976; // @[TLSimpleL2.scala 586:43:freechips.rocketchip.system.DefaultConfig.fir@224790.4]
  assign _T_14172 = _T_274 & _T_14180; // @[TLSimpleL2.scala 590:54:freechips.rocketchip.system.DefaultConfig.fir@224794.4]
  assign _T_14174 = value_2 == 3'h7; // @[Counter.scala 34:24:freechips.rocketchip.system.DefaultConfig.fir@224797.6]
  assign _T_14176 = value_2 + 3'h1; // @[Counter.scala 35:22:freechips.rocketchip.system.DefaultConfig.fir@224799.6]
  assign _T_14177 = _T_14172 & _T_14174; // @[Counter.scala 64:20:freechips.rocketchip.system.DefaultConfig.fir@224802.4]
  assign _T_14179 = _T_14180 & _T_14177; // @[TLSimpleL2.scala 591:38:freechips.rocketchip.system.DefaultConfig.fir@224804.4]
  assign _GEN_6979 = _T_14179 ? 4'hc : _GEN_6977; // @[TLSimpleL2.scala 591:50:freechips.rocketchip.system.DefaultConfig.fir@224805.4]
  assign _T_14182 = _T_14269 & _T_14168; // @[TLSimpleL2.scala 597:40:freechips.rocketchip.system.DefaultConfig.fir@224810.4]
  assign _T_14188 = _T_14199 & _T_274; // @[TLSimpleL2.scala 612:42:freechips.rocketchip.system.DefaultConfig.fir@224827.4]
  assign _T_14190 = _T_14168 & _T_14268; // @[TLSimpleL2.scala 615:62:freechips.rocketchip.system.DefaultConfig.fir@224832.4]
  assign _T_14192 = value_3 == 3'h7; // @[Counter.scala 34:24:freechips.rocketchip.system.DefaultConfig.fir@224835.6]
  assign _T_14194 = value_3 + 3'h1; // @[Counter.scala 35:22:freechips.rocketchip.system.DefaultConfig.fir@224837.6]
  assign _T_14195 = _T_14190 & _T_14192; // @[Counter.scala 64:20:freechips.rocketchip.system.DefaultConfig.fir@224840.4]
  assign _T_14197 = _T_14268 & _T_14168; // @[TLSimpleL2.scala 616:37:freechips.rocketchip.system.DefaultConfig.fir@224842.4]
  assign _GEN_7004 = 3'h1 == value_2 ? _T_14075_1 : _T_14075_0; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  assign _GEN_7005 = 3'h2 == value_2 ? _T_14075_2 : _GEN_7004; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  assign _GEN_7006 = 3'h3 == value_2 ? _T_14075_3 : _GEN_7005; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  assign _GEN_7007 = 3'h4 == value_2 ? _T_14075_4 : _GEN_7006; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  assign _GEN_7008 = 3'h5 == value_2 ? _T_14075_5 : _GEN_7007; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  assign _GEN_7009 = 3'h6 == value_2 ? _T_14075_6 : _GEN_7008; // @[TLSimpleL2.scala 640:26:freechips.rocketchip.system.DefaultConfig.fir@224928.4]
  assign _T_14272 = _T_14286 & _T_289; // @[TLSimpleL2.scala 652:35:freechips.rocketchip.system.DefaultConfig.fir@224937.4]
  assign _T_14274 = _T_320 + 3'h1; // @[TLSimpleL2.scala 653:42:freechips.rocketchip.system.DefaultConfig.fir@224940.6]
  assign _T_14283 = {{1'd0}, _T_320}; // @[TLSimpleL2.scala 661:64:freechips.rocketchip.system.DefaultConfig.fir@224949.4]
  assign _T_14284 = _T_14283[2:0]; // @[TLSimpleL2.scala 661:64:freechips.rocketchip.system.DefaultConfig.fir@224950.4]
  assign _GEN_7015 = 3'h1 == _T_14284 ? _T_14075_1 : _T_14075_0; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  assign _GEN_7016 = 3'h2 == _T_14284 ? _T_14075_2 : _GEN_7015; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  assign _GEN_7017 = 3'h3 == _T_14284 ? _T_14075_3 : _GEN_7016; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  assign _GEN_7018 = 3'h4 == _T_14284 ? _T_14075_4 : _GEN_7017; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  assign _GEN_7019 = 3'h5 == _T_14284 ? _T_14075_5 : _GEN_7018; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  assign _GEN_7020 = 3'h6 == _T_14284 ? _T_14075_6 : _GEN_7019; // @[TLSimpleL2.scala 661:22:freechips.rocketchip.system.DefaultConfig.fir@224951.4]
  assign auto_in_a_ready = _T_451 | _T_426; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultConfig.fir@221007.4]
  assign auto_in_d_valid = _T_456 | _T_14286; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultConfig.fir@221007.4]
  assign auto_in_d_bits_opcode = {{2'd0}, _T_14286}; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultConfig.fir@221007.4]
  assign auto_in_d_bits_size = _T_299; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultConfig.fir@221007.4]
  assign auto_in_d_bits_source = _T_293; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultConfig.fir@221007.4]
  assign auto_in_d_bits_data = 3'h7 == _T_14284 ? _T_14075_7 : _GEN_7020; // @[LazyModule.scala 173:31:freechips.rocketchip.system.DefaultConfig.fir@221007.4]
  assign auto_out_a_valid = _T_14180 | _T_14199; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultConfig.fir@221006.4]
  assign auto_out_a_bits_opcode = _T_14199 ? 3'h4 : 3'h0; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultConfig.fir@221006.4]
  assign auto_out_a_bits_address = _T_14199 ? _T_14164 : _T_13374; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultConfig.fir@221006.4]
  assign auto_out_a_bits_data = 3'h7 == value_2 ? _T_14075_7 : _GEN_7009; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultConfig.fir@221006.4]
  assign auto_out_d_ready = _T_14268 | _T_14269; // @[LazyModule.scala 173:49:freechips.rocketchip.system.DefaultConfig.fir@221006.4]
  assign cp_capacity = 4'hf == cp_capacity_dsid ? _T_13304_15 : _GEN_6289; // @[TLSimpleL2.scala 361:19:freechips.rocketchip.system.DefaultConfig.fir@223687.4]
  assign TLMonitor_clock = clock; // @[:freechips.rocketchip.system.DefaultConfig.fir@220969.4]
  assign TLMonitor_reset = reset; // @[:freechips.rocketchip.system.DefaultConfig.fir@220970.4]
  assign TLMonitor_io_in_a_ready = _T_451 | _T_426; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_valid = auto_in_a_valid; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_opcode = auto_in_a_bits_opcode; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_param = auto_in_a_bits_param; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_size = auto_in_a_bits_size; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_source = auto_in_a_bits_source; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_address = auto_in_a_bits_address; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_mask = auto_in_a_bits_mask; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_a_bits_corrupt = auto_in_a_bits_corrupt; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_d_ready = auto_in_d_ready; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_d_valid = _T_456 | _T_14286; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_d_bits_opcode = {{2'd0}, _T_14286}; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_d_bits_size = _T_299; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign TLMonitor_io_in_d_bits_source = _T_293; // @[Nodes.scala 26:19:freechips.rocketchip.system.DefaultConfig.fir@221003.4]
  assign L2_meta_array_RW0_wdata_0_valid = _T_262 ? 1'h0 : _GEN_6312; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_0_dirty = _T_262 ? 1'h0 : _GEN_6313; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_0_tag = _T_262 ? 16'h0 : _GEN_6314; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_0_rr_state = _T_262 ? 1'h0 : _T_13461; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_0_dsid = _T_13584_0_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_1_valid = _T_262 ? 1'h0 : _GEN_6316; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_1_dirty = _T_262 ? 1'h0 : _GEN_6317; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_1_tag = _T_262 ? 16'h0 : _GEN_6318; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_1_rr_state = _T_262 ? 1'h0 : _T_13469; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_1_dsid = _T_13584_1_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_2_valid = _T_262 ? 1'h0 : _GEN_6320; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_2_dirty = _T_262 ? 1'h0 : _GEN_6321; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_2_tag = _T_262 ? 16'h0 : _GEN_6322; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_2_rr_state = _T_262 ? 1'h0 : _T_13477; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_2_dsid = _T_13584_2_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_3_valid = _T_262 ? 1'h0 : _GEN_6324; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_3_dirty = _T_262 ? 1'h0 : _GEN_6325; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_3_tag = _T_262 ? 16'h0 : _GEN_6326; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_3_rr_state = _T_262 ? 1'h0 : _T_13485; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_3_dsid = _T_13584_3_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_4_valid = _T_262 ? 1'h0 : _GEN_6328; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_4_dirty = _T_262 ? 1'h0 : _GEN_6329; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_4_tag = _T_262 ? 16'h0 : _GEN_6330; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_4_rr_state = _T_262 ? 1'h0 : _T_13493; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_4_dsid = _T_13584_4_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_5_valid = _T_262 ? 1'h0 : _GEN_6332; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_5_dirty = _T_262 ? 1'h0 : _GEN_6333; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_5_tag = _T_262 ? 16'h0 : _GEN_6334; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_5_rr_state = _T_262 ? 1'h0 : _T_13501; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_5_dsid = _T_13584_5_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_6_valid = _T_262 ? 1'h0 : _GEN_6336; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_6_dirty = _T_262 ? 1'h0 : _GEN_6337; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_6_tag = _T_262 ? 16'h0 : _GEN_6338; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_6_rr_state = _T_262 ? 1'h0 : _T_13509; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_6_dsid = _T_13584_6_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_7_valid = _T_262 ? 1'h0 : _GEN_6340; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_7_dirty = _T_262 ? 1'h0 : _GEN_6341; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_7_tag = _T_262 ? 16'h0 : _GEN_6342; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_7_rr_state = _T_262 ? 1'h0 : _T_13517; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_7_dsid = _T_13584_7_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_8_valid = _T_262 ? 1'h0 : _GEN_6344; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_8_dirty = _T_262 ? 1'h0 : _GEN_6345; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_8_tag = _T_262 ? 16'h0 : _GEN_6346; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_8_rr_state = _T_262 ? 1'h0 : _T_13525; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_8_dsid = _T_13584_8_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_9_valid = _T_262 ? 1'h0 : _GEN_6348; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_9_dirty = _T_262 ? 1'h0 : _GEN_6349; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_9_tag = _T_262 ? 16'h0 : _GEN_6350; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_9_rr_state = _T_262 ? 1'h0 : _T_13533; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_9_dsid = _T_13584_9_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_10_valid = _T_262 ? 1'h0 : _GEN_6352; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_10_dirty = _T_262 ? 1'h0 : _GEN_6353; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_10_tag = _T_262 ? 16'h0 : _GEN_6354; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_10_rr_state = _T_262 ? 1'h0 : _T_13541; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_10_dsid = _T_13584_10_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_11_valid = _T_262 ? 1'h0 : _GEN_6356; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_11_dirty = _T_262 ? 1'h0 : _GEN_6357; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_11_tag = _T_262 ? 16'h0 : _GEN_6358; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_11_rr_state = _T_262 ? 1'h0 : _T_13549; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_11_dsid = _T_13584_11_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_12_valid = _T_262 ? 1'h0 : _GEN_6360; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_12_dirty = _T_262 ? 1'h0 : _GEN_6361; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_12_tag = _T_262 ? 16'h0 : _GEN_6362; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_12_rr_state = _T_262 ? 1'h0 : _T_13557; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_12_dsid = _T_13584_12_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_13_valid = _T_262 ? 1'h0 : _GEN_6364; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_13_dirty = _T_262 ? 1'h0 : _GEN_6365; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_13_tag = _T_262 ? 16'h0 : _GEN_6366; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_13_rr_state = _T_262 ? 1'h0 : _T_13565; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_13_dsid = _T_13584_13_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_14_valid = _T_262 ? 1'h0 : _GEN_6368; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_14_dirty = _T_262 ? 1'h0 : _GEN_6369; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_14_tag = _T_262 ? 16'h0 : _GEN_6370; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_14_rr_state = _T_262 ? 1'h0 : _T_13573; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_14_dsid = _T_13584_14_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_15_valid = _T_262 ? 1'h0 : _GEN_6372; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_15_dirty = _T_262 ? 1'h0 : _GEN_6373; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_15_tag = _T_262 ? 16'h0 : _GEN_6374; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_15_rr_state = _T_262 ? 1'h0 : _T_13581; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_meta_array_RW0_wdata_15_dsid = _T_13584_15_dsid[3:0]; // @[:freechips.rocketchip.system.DefaultConfig.fir@224180.6]
  assign L2_data_array_RW0_wdata_0 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224596.8]
  assign L2_data_array_RW0_wdata_1 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224599.8]
  assign L2_data_array_RW0_wdata_2 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224602.8]
  assign L2_data_array_RW0_wdata_3 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224605.8]
  assign L2_data_array_RW0_wdata_4 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224608.8]
  assign L2_data_array_RW0_wdata_5 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224611.8]
  assign L2_data_array_RW0_wdata_6 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224614.8]
  assign L2_data_array_RW0_wdata_7 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224617.8]
  assign L2_data_array_RW0_wdata_8 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224620.8]
  assign L2_data_array_RW0_wdata_9 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224623.8]
  assign L2_data_array_RW0_wdata_10 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224626.8]
  assign L2_data_array_RW0_wdata_11 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224629.8]
  assign L2_data_array_RW0_wdata_12 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224632.8]
  assign L2_data_array_RW0_wdata_13 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224635.8]
  assign L2_data_array_RW0_wdata_14 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224638.8]
  assign L2_data_array_RW0_wdata_15 = 3'h7 == _T_14157 ? _T_14075_7 : _GEN_6973; // @[:freechips.rocketchip.system.DefaultConfig.fir@224641.8]
  assign L2_data_array_RW0_wmask_0 = _T_13909 == 4'h0; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224596.8]
  assign L2_data_array_RW0_wmask_1 = _T_13909 == 4'h1; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224599.8]
  assign L2_data_array_RW0_wmask_2 = _T_13909 == 4'h2; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224602.8]
  assign L2_data_array_RW0_wmask_3 = _T_13909 == 4'h3; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224605.8]
  assign L2_data_array_RW0_wmask_4 = _T_13909 == 4'h4; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224608.8]
  assign L2_data_array_RW0_wmask_5 = _T_13909 == 4'h5; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224611.8]
  assign L2_data_array_RW0_wmask_6 = _T_13909 == 4'h6; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224614.8]
  assign L2_data_array_RW0_wmask_7 = _T_13909 == 4'h7; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224617.8]
  assign L2_data_array_RW0_wmask_8 = _T_13909 == 4'h8; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224620.8]
  assign L2_data_array_RW0_wmask_9 = _T_13909 == 4'h9; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224623.8]
  assign L2_data_array_RW0_wmask_10 = _T_13909 == 4'ha; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224626.8]
  assign L2_data_array_RW0_wmask_11 = _T_13909 == 4'hb; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224629.8]
  assign L2_data_array_RW0_wmask_12 = _T_13909 == 4'hc; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224632.8]
  assign L2_data_array_RW0_wmask_13 = _T_13909 == 4'hd; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224635.8]
  assign L2_data_array_RW0_wmask_14 = _T_13909 == 4'he; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224638.8]
  assign L2_data_array_RW0_wmask_15 = _T_13909 == 4'hf; // @[:freechips.rocketchip.system.DefaultConfig.fir@224594.6 :freechips.rocketchip.system.DefaultConfig.fir@224641.8]
  assign _GEN_7033 = _T_335 == 1'h0; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  assign _GEN_7034 = _T_429 & _GEN_7033; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  assign _GEN_7035 = _T_426 == 1'h0; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  assign _GEN_7036 = _GEN_7034 & _GEN_7035; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
  assign _GEN_7041 = _T_13383 == 1'h0; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  assign _GEN_7042 = _T_482 & _GEN_7041; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  assign _GEN_7043 = _T_13392 == 1'h0; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  assign _GEN_7044 = _GEN_7042 & _GEN_7043; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
  assign _GEN_7049 = _T_483 & _T_13659; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224190.10]
  assign _GEN_7051 = _T_13896 & _T_14097; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7052 = _T_13153 == 1'h0; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7053 = _GEN_7051 & _GEN_7052; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7054 = _T_14098 == 1'h0; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7055 = _GEN_7053 & _GEN_7054; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7056 = _T_13154 == 1'h0; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7057 = _GEN_7055 & _GEN_7056; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
  assign _GEN_7066 = _T_14182 & _GEN_7054; // @[TLSimpleL2.scala 602:17:freechips.rocketchip.system.DefaultConfig.fir@224821.10]
  assign L2_meta_array_RW0_wmode = _T_262 | _T_482;
  assign L2_meta_array_RW0_clk = clock;
  assign L2_meta_array_RW0_en = _T_486 | _T_483;
  assign L2_meta_array_RW0_addr = _T_483 ? _T_13620 : _T_481;
  assign L2_data_array_RW0_wmode = _T_267 == 4'h9;
  assign L2_data_array_RW0_clk = clock;
  assign L2_data_array_RW0_en = _T_14021 | _T_13912;
  assign L2_data_array_RW0_addr = _T_13912 ? _T_13914 : _T_13901;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_258 = _RAND_0[12:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_267 = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {2{`RANDOM}};
  _T_291 = _RAND_2[32:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  _T_293 = _RAND_3[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  _T_297 = _RAND_4[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  _T_299 = _RAND_5[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_301 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_303 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  _T_306 = _RAND_8[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  _T_312 = _RAND_9[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  _T_317 = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  _T_320 = _RAND_11[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {2{`RANDOM}};
  _T_344_0 = _RAND_12[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_344_1 = _RAND_13[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {2{`RANDOM}};
  _T_344_2 = _RAND_14[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_344_3 = _RAND_15[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_344_4 = _RAND_16[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_344_5 = _RAND_17[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_344_6 = _RAND_18[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_344_7 = _RAND_19[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_397_0 = _RAND_20[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_397_1 = _RAND_21[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  _T_397_2 = _RAND_22[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  _T_397_3 = _RAND_23[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  _T_397_4 = _RAND_24[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  _T_397_5 = _RAND_25[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  _T_397_6 = _RAND_26[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  _T_397_7 = _RAND_27[7:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  _T_684 = _RAND_28[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  _T_686 = _RAND_29[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  _T_690_0 = _RAND_30[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  _T_690_1 = _RAND_31[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  _T_690_2 = _RAND_32[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  _T_690_3 = _RAND_33[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  _T_690_4 = _RAND_34[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  _T_690_5 = _RAND_35[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  _T_690_6 = _RAND_36[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_690_7 = _RAND_37[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_690_8 = _RAND_38[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_690_9 = _RAND_39[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_690_10 = _RAND_40[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_690_11 = _RAND_41[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_690_12 = _RAND_42[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  _T_690_13 = _RAND_43[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  _T_690_14 = _RAND_44[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  _T_690_15 = _RAND_45[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  _T_710 = _RAND_46[15:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  _T_714_0 = _RAND_47[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  _T_714_1 = _RAND_48[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  _T_714_2 = _RAND_49[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  _T_714_3 = _RAND_50[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  _T_714_4 = _RAND_51[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  _T_714_5 = _RAND_52[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  _T_714_6 = _RAND_53[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  _T_714_7 = _RAND_54[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  _T_714_8 = _RAND_55[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  _T_714_9 = _RAND_56[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  _T_714_10 = _RAND_57[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  _T_714_11 = _RAND_58[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  _T_714_12 = _RAND_59[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  _T_714_13 = _RAND_60[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  _T_714_14 = _RAND_61[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  _T_714_15 = _RAND_62[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  _T_6887_0 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  _T_6887_1 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  _T_6887_2 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  _T_6887_3 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  _T_6887_4 = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  _T_6887_5 = _RAND_68[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  _T_6887_6 = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  _T_6887_7 = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  _T_6887_8 = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  _T_6887_9 = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_6887_10 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_6887_11 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_6887_12 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_6887_13 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_6887_14 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  _T_6887_15 = _RAND_78[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  _T_6887_16 = _RAND_79[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  _T_6887_17 = _RAND_80[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  _T_6887_18 = _RAND_81[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  _T_6887_19 = _RAND_82[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  _T_6887_20 = _RAND_83[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  _T_6887_21 = _RAND_84[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  _T_6887_22 = _RAND_85[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  _T_6887_23 = _RAND_86[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  _T_6887_24 = _RAND_87[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  _T_6887_25 = _RAND_88[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  _T_6887_26 = _RAND_89[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  _T_6887_27 = _RAND_90[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  _T_6887_28 = _RAND_91[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  _T_6887_29 = _RAND_92[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  _T_6887_30 = _RAND_93[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  _T_6887_31 = _RAND_94[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  _T_6887_32 = _RAND_95[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  _T_6887_33 = _RAND_96[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  _T_6887_34 = _RAND_97[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  _T_6887_35 = _RAND_98[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  _T_6887_36 = _RAND_99[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  _T_6887_37 = _RAND_100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  _T_6887_38 = _RAND_101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  _T_6887_39 = _RAND_102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  _T_6887_40 = _RAND_103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  _T_6887_41 = _RAND_104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  _T_6887_42 = _RAND_105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  _T_6887_43 = _RAND_106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  _T_6887_44 = _RAND_107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  _T_6887_45 = _RAND_108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  _T_6887_46 = _RAND_109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  _T_6887_47 = _RAND_110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  _T_6887_48 = _RAND_111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  _T_6887_49 = _RAND_112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  _T_6887_50 = _RAND_113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  _T_6887_51 = _RAND_114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  _T_6887_52 = _RAND_115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  _T_6887_53 = _RAND_116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  _T_6887_54 = _RAND_117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  _T_6887_55 = _RAND_118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  _T_6887_56 = _RAND_119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  _T_6887_57 = _RAND_120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  _T_6887_58 = _RAND_121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  _T_6887_59 = _RAND_122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  _T_6887_60 = _RAND_123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  _T_6887_61 = _RAND_124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  _T_6887_62 = _RAND_125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  _T_6887_63 = _RAND_126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  _T_6887_64 = _RAND_127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  _T_6887_65 = _RAND_128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  _T_6887_66 = _RAND_129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  _T_6887_67 = _RAND_130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  _T_6887_68 = _RAND_131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  _T_6887_69 = _RAND_132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  _T_6887_70 = _RAND_133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  _T_6887_71 = _RAND_134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  _T_6887_72 = _RAND_135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  _T_6887_73 = _RAND_136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  _T_6887_74 = _RAND_137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  _T_6887_75 = _RAND_138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  _T_6887_76 = _RAND_139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  _T_6887_77 = _RAND_140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  _T_6887_78 = _RAND_141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  _T_6887_79 = _RAND_142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  _T_6887_80 = _RAND_143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  _T_6887_81 = _RAND_144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  _T_6887_82 = _RAND_145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  _T_6887_83 = _RAND_146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  _T_6887_84 = _RAND_147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  _T_6887_85 = _RAND_148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  _T_6887_86 = _RAND_149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  _T_6887_87 = _RAND_150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  _T_6887_88 = _RAND_151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  _T_6887_89 = _RAND_152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  _T_6887_90 = _RAND_153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  _T_6887_91 = _RAND_154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  _T_6887_92 = _RAND_155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  _T_6887_93 = _RAND_156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  _T_6887_94 = _RAND_157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  _T_6887_95 = _RAND_158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  _T_6887_96 = _RAND_159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  _T_6887_97 = _RAND_160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  _T_6887_98 = _RAND_161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  _T_6887_99 = _RAND_162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  _T_6887_100 = _RAND_163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  _T_6887_101 = _RAND_164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  _T_6887_102 = _RAND_165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  _T_6887_103 = _RAND_166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  _T_6887_104 = _RAND_167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  _T_6887_105 = _RAND_168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  _T_6887_106 = _RAND_169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  _T_6887_107 = _RAND_170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  _T_6887_108 = _RAND_171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  _T_6887_109 = _RAND_172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  _T_6887_110 = _RAND_173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  _T_6887_111 = _RAND_174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  _T_6887_112 = _RAND_175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  _T_6887_113 = _RAND_176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  _T_6887_114 = _RAND_177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  _T_6887_115 = _RAND_178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  _T_6887_116 = _RAND_179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  _T_6887_117 = _RAND_180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  _T_6887_118 = _RAND_181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  _T_6887_119 = _RAND_182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  _T_6887_120 = _RAND_183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  _T_6887_121 = _RAND_184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  _T_6887_122 = _RAND_185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  _T_6887_123 = _RAND_186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  _T_6887_124 = _RAND_187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  _T_6887_125 = _RAND_188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  _T_6887_126 = _RAND_189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  _T_6887_127 = _RAND_190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  _T_6887_128 = _RAND_191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  _T_6887_129 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  _T_6887_130 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  _T_6887_131 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  _T_6887_132 = _RAND_195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  _T_6887_133 = _RAND_196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  _T_6887_134 = _RAND_197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  _T_6887_135 = _RAND_198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  _T_6887_136 = _RAND_199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  _T_6887_137 = _RAND_200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  _T_6887_138 = _RAND_201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  _T_6887_139 = _RAND_202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  _T_6887_140 = _RAND_203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  _T_6887_141 = _RAND_204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  _T_6887_142 = _RAND_205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  _T_6887_143 = _RAND_206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  _T_6887_144 = _RAND_207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  _T_6887_145 = _RAND_208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  _T_6887_146 = _RAND_209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  _T_6887_147 = _RAND_210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  _T_6887_148 = _RAND_211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  _T_6887_149 = _RAND_212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  _T_6887_150 = _RAND_213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  _T_6887_151 = _RAND_214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  _T_6887_152 = _RAND_215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  _T_6887_153 = _RAND_216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  _T_6887_154 = _RAND_217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  _T_6887_155 = _RAND_218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  _T_6887_156 = _RAND_219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  _T_6887_157 = _RAND_220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  _T_6887_158 = _RAND_221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  _T_6887_159 = _RAND_222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  _T_6887_160 = _RAND_223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  _T_6887_161 = _RAND_224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  _T_6887_162 = _RAND_225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  _T_6887_163 = _RAND_226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  _T_6887_164 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  _T_6887_165 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  _T_6887_166 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  _T_6887_167 = _RAND_230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  _T_6887_168 = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  _T_6887_169 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  _T_6887_170 = _RAND_233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  _T_6887_171 = _RAND_234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  _T_6887_172 = _RAND_235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  _T_6887_173 = _RAND_236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  _T_6887_174 = _RAND_237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  _T_6887_175 = _RAND_238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  _T_6887_176 = _RAND_239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  _T_6887_177 = _RAND_240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  _T_6887_178 = _RAND_241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  _T_6887_179 = _RAND_242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  _T_6887_180 = _RAND_243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  _T_6887_181 = _RAND_244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  _T_6887_182 = _RAND_245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  _T_6887_183 = _RAND_246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  _T_6887_184 = _RAND_247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  _T_6887_185 = _RAND_248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  _T_6887_186 = _RAND_249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  _T_6887_187 = _RAND_250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  _T_6887_188 = _RAND_251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  _T_6887_189 = _RAND_252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  _T_6887_190 = _RAND_253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  _T_6887_191 = _RAND_254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  _T_6887_192 = _RAND_255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  _T_6887_193 = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  _T_6887_194 = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  _T_6887_195 = _RAND_258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  _T_6887_196 = _RAND_259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  _T_6887_197 = _RAND_260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  _T_6887_198 = _RAND_261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  _T_6887_199 = _RAND_262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  _T_6887_200 = _RAND_263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  _T_6887_201 = _RAND_264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  _T_6887_202 = _RAND_265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  _T_6887_203 = _RAND_266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  _T_6887_204 = _RAND_267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  _T_6887_205 = _RAND_268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  _T_6887_206 = _RAND_269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  _T_6887_207 = _RAND_270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  _T_6887_208 = _RAND_271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  _T_6887_209 = _RAND_272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  _T_6887_210 = _RAND_273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  _T_6887_211 = _RAND_274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  _T_6887_212 = _RAND_275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  _T_6887_213 = _RAND_276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  _T_6887_214 = _RAND_277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  _T_6887_215 = _RAND_278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  _T_6887_216 = _RAND_279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  _T_6887_217 = _RAND_280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  _T_6887_218 = _RAND_281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  _T_6887_219 = _RAND_282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  _T_6887_220 = _RAND_283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  _T_6887_221 = _RAND_284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  _T_6887_222 = _RAND_285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  _T_6887_223 = _RAND_286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  _T_6887_224 = _RAND_287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  _T_6887_225 = _RAND_288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  _T_6887_226 = _RAND_289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  _T_6887_227 = _RAND_290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  _T_6887_228 = _RAND_291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  _T_6887_229 = _RAND_292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  _T_6887_230 = _RAND_293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  _T_6887_231 = _RAND_294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  _T_6887_232 = _RAND_295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  _T_6887_233 = _RAND_296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  _T_6887_234 = _RAND_297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  _T_6887_235 = _RAND_298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  _T_6887_236 = _RAND_299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  _T_6887_237 = _RAND_300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  _T_6887_238 = _RAND_301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  _T_6887_239 = _RAND_302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  _T_6887_240 = _RAND_303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  _T_6887_241 = _RAND_304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  _T_6887_242 = _RAND_305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  _T_6887_243 = _RAND_306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  _T_6887_244 = _RAND_307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  _T_6887_245 = _RAND_308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  _T_6887_246 = _RAND_309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  _T_6887_247 = _RAND_310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  _T_6887_248 = _RAND_311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  _T_6887_249 = _RAND_312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  _T_6887_250 = _RAND_313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  _T_6887_251 = _RAND_314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  _T_6887_252 = _RAND_315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  _T_6887_253 = _RAND_316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  _T_6887_254 = _RAND_317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  _T_6887_255 = _RAND_318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  _T_6887_256 = _RAND_319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  _T_6887_257 = _RAND_320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  _T_6887_258 = _RAND_321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  _T_6887_259 = _RAND_322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  _T_6887_260 = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  _T_6887_261 = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  _T_6887_262 = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  _T_6887_263 = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  _T_6887_264 = _RAND_327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  _T_6887_265 = _RAND_328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  _T_6887_266 = _RAND_329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  _T_6887_267 = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  _T_6887_268 = _RAND_331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  _T_6887_269 = _RAND_332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_333 = {1{`RANDOM}};
  _T_6887_270 = _RAND_333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_334 = {1{`RANDOM}};
  _T_6887_271 = _RAND_334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_335 = {1{`RANDOM}};
  _T_6887_272 = _RAND_335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_336 = {1{`RANDOM}};
  _T_6887_273 = _RAND_336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_337 = {1{`RANDOM}};
  _T_6887_274 = _RAND_337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_338 = {1{`RANDOM}};
  _T_6887_275 = _RAND_338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_339 = {1{`RANDOM}};
  _T_6887_276 = _RAND_339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_340 = {1{`RANDOM}};
  _T_6887_277 = _RAND_340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_341 = {1{`RANDOM}};
  _T_6887_278 = _RAND_341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_342 = {1{`RANDOM}};
  _T_6887_279 = _RAND_342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_343 = {1{`RANDOM}};
  _T_6887_280 = _RAND_343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_344 = {1{`RANDOM}};
  _T_6887_281 = _RAND_344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_345 = {1{`RANDOM}};
  _T_6887_282 = _RAND_345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_346 = {1{`RANDOM}};
  _T_6887_283 = _RAND_346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_347 = {1{`RANDOM}};
  _T_6887_284 = _RAND_347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_348 = {1{`RANDOM}};
  _T_6887_285 = _RAND_348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_349 = {1{`RANDOM}};
  _T_6887_286 = _RAND_349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_350 = {1{`RANDOM}};
  _T_6887_287 = _RAND_350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_351 = {1{`RANDOM}};
  _T_6887_288 = _RAND_351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_352 = {1{`RANDOM}};
  _T_6887_289 = _RAND_352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_353 = {1{`RANDOM}};
  _T_6887_290 = _RAND_353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_354 = {1{`RANDOM}};
  _T_6887_291 = _RAND_354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_355 = {1{`RANDOM}};
  _T_6887_292 = _RAND_355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_356 = {1{`RANDOM}};
  _T_6887_293 = _RAND_356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_357 = {1{`RANDOM}};
  _T_6887_294 = _RAND_357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_358 = {1{`RANDOM}};
  _T_6887_295 = _RAND_358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_359 = {1{`RANDOM}};
  _T_6887_296 = _RAND_359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_360 = {1{`RANDOM}};
  _T_6887_297 = _RAND_360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_361 = {1{`RANDOM}};
  _T_6887_298 = _RAND_361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_362 = {1{`RANDOM}};
  _T_6887_299 = _RAND_362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_363 = {1{`RANDOM}};
  _T_6887_300 = _RAND_363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_364 = {1{`RANDOM}};
  _T_6887_301 = _RAND_364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_365 = {1{`RANDOM}};
  _T_6887_302 = _RAND_365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_366 = {1{`RANDOM}};
  _T_6887_303 = _RAND_366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_367 = {1{`RANDOM}};
  _T_6887_304 = _RAND_367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_368 = {1{`RANDOM}};
  _T_6887_305 = _RAND_368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_369 = {1{`RANDOM}};
  _T_6887_306 = _RAND_369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_370 = {1{`RANDOM}};
  _T_6887_307 = _RAND_370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_371 = {1{`RANDOM}};
  _T_6887_308 = _RAND_371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_372 = {1{`RANDOM}};
  _T_6887_309 = _RAND_372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_373 = {1{`RANDOM}};
  _T_6887_310 = _RAND_373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_374 = {1{`RANDOM}};
  _T_6887_311 = _RAND_374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_375 = {1{`RANDOM}};
  _T_6887_312 = _RAND_375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_376 = {1{`RANDOM}};
  _T_6887_313 = _RAND_376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_377 = {1{`RANDOM}};
  _T_6887_314 = _RAND_377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_378 = {1{`RANDOM}};
  _T_6887_315 = _RAND_378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_379 = {1{`RANDOM}};
  _T_6887_316 = _RAND_379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_380 = {1{`RANDOM}};
  _T_6887_317 = _RAND_380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_381 = {1{`RANDOM}};
  _T_6887_318 = _RAND_381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_382 = {1{`RANDOM}};
  _T_6887_319 = _RAND_382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_383 = {1{`RANDOM}};
  _T_6887_320 = _RAND_383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_384 = {1{`RANDOM}};
  _T_6887_321 = _RAND_384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_385 = {1{`RANDOM}};
  _T_6887_322 = _RAND_385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_386 = {1{`RANDOM}};
  _T_6887_323 = _RAND_386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_387 = {1{`RANDOM}};
  _T_6887_324 = _RAND_387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_388 = {1{`RANDOM}};
  _T_6887_325 = _RAND_388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_389 = {1{`RANDOM}};
  _T_6887_326 = _RAND_389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_390 = {1{`RANDOM}};
  _T_6887_327 = _RAND_390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_391 = {1{`RANDOM}};
  _T_6887_328 = _RAND_391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_392 = {1{`RANDOM}};
  _T_6887_329 = _RAND_392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_393 = {1{`RANDOM}};
  _T_6887_330 = _RAND_393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_394 = {1{`RANDOM}};
  _T_6887_331 = _RAND_394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_395 = {1{`RANDOM}};
  _T_6887_332 = _RAND_395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_396 = {1{`RANDOM}};
  _T_6887_333 = _RAND_396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_397 = {1{`RANDOM}};
  _T_6887_334 = _RAND_397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_398 = {1{`RANDOM}};
  _T_6887_335 = _RAND_398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_399 = {1{`RANDOM}};
  _T_6887_336 = _RAND_399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_400 = {1{`RANDOM}};
  _T_6887_337 = _RAND_400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_401 = {1{`RANDOM}};
  _T_6887_338 = _RAND_401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_402 = {1{`RANDOM}};
  _T_6887_339 = _RAND_402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_403 = {1{`RANDOM}};
  _T_6887_340 = _RAND_403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_404 = {1{`RANDOM}};
  _T_6887_341 = _RAND_404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_405 = {1{`RANDOM}};
  _T_6887_342 = _RAND_405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_406 = {1{`RANDOM}};
  _T_6887_343 = _RAND_406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_407 = {1{`RANDOM}};
  _T_6887_344 = _RAND_407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_408 = {1{`RANDOM}};
  _T_6887_345 = _RAND_408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_409 = {1{`RANDOM}};
  _T_6887_346 = _RAND_409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_410 = {1{`RANDOM}};
  _T_6887_347 = _RAND_410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_411 = {1{`RANDOM}};
  _T_6887_348 = _RAND_411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_412 = {1{`RANDOM}};
  _T_6887_349 = _RAND_412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_413 = {1{`RANDOM}};
  _T_6887_350 = _RAND_413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_414 = {1{`RANDOM}};
  _T_6887_351 = _RAND_414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_415 = {1{`RANDOM}};
  _T_6887_352 = _RAND_415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_416 = {1{`RANDOM}};
  _T_6887_353 = _RAND_416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_417 = {1{`RANDOM}};
  _T_6887_354 = _RAND_417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_418 = {1{`RANDOM}};
  _T_6887_355 = _RAND_418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_419 = {1{`RANDOM}};
  _T_6887_356 = _RAND_419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_420 = {1{`RANDOM}};
  _T_6887_357 = _RAND_420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_421 = {1{`RANDOM}};
  _T_6887_358 = _RAND_421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_422 = {1{`RANDOM}};
  _T_6887_359 = _RAND_422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_423 = {1{`RANDOM}};
  _T_6887_360 = _RAND_423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_424 = {1{`RANDOM}};
  _T_6887_361 = _RAND_424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_425 = {1{`RANDOM}};
  _T_6887_362 = _RAND_425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_426 = {1{`RANDOM}};
  _T_6887_363 = _RAND_426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_427 = {1{`RANDOM}};
  _T_6887_364 = _RAND_427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_428 = {1{`RANDOM}};
  _T_6887_365 = _RAND_428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_429 = {1{`RANDOM}};
  _T_6887_366 = _RAND_429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_430 = {1{`RANDOM}};
  _T_6887_367 = _RAND_430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_431 = {1{`RANDOM}};
  _T_6887_368 = _RAND_431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_432 = {1{`RANDOM}};
  _T_6887_369 = _RAND_432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_433 = {1{`RANDOM}};
  _T_6887_370 = _RAND_433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_434 = {1{`RANDOM}};
  _T_6887_371 = _RAND_434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_435 = {1{`RANDOM}};
  _T_6887_372 = _RAND_435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_436 = {1{`RANDOM}};
  _T_6887_373 = _RAND_436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_437 = {1{`RANDOM}};
  _T_6887_374 = _RAND_437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_438 = {1{`RANDOM}};
  _T_6887_375 = _RAND_438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_439 = {1{`RANDOM}};
  _T_6887_376 = _RAND_439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_440 = {1{`RANDOM}};
  _T_6887_377 = _RAND_440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_441 = {1{`RANDOM}};
  _T_6887_378 = _RAND_441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_442 = {1{`RANDOM}};
  _T_6887_379 = _RAND_442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_443 = {1{`RANDOM}};
  _T_6887_380 = _RAND_443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_444 = {1{`RANDOM}};
  _T_6887_381 = _RAND_444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_445 = {1{`RANDOM}};
  _T_6887_382 = _RAND_445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_446 = {1{`RANDOM}};
  _T_6887_383 = _RAND_446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_447 = {1{`RANDOM}};
  _T_6887_384 = _RAND_447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_448 = {1{`RANDOM}};
  _T_6887_385 = _RAND_448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_449 = {1{`RANDOM}};
  _T_6887_386 = _RAND_449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_450 = {1{`RANDOM}};
  _T_6887_387 = _RAND_450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_451 = {1{`RANDOM}};
  _T_6887_388 = _RAND_451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_452 = {1{`RANDOM}};
  _T_6887_389 = _RAND_452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_453 = {1{`RANDOM}};
  _T_6887_390 = _RAND_453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_454 = {1{`RANDOM}};
  _T_6887_391 = _RAND_454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_455 = {1{`RANDOM}};
  _T_6887_392 = _RAND_455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_456 = {1{`RANDOM}};
  _T_6887_393 = _RAND_456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_457 = {1{`RANDOM}};
  _T_6887_394 = _RAND_457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_458 = {1{`RANDOM}};
  _T_6887_395 = _RAND_458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_459 = {1{`RANDOM}};
  _T_6887_396 = _RAND_459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_460 = {1{`RANDOM}};
  _T_6887_397 = _RAND_460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_461 = {1{`RANDOM}};
  _T_6887_398 = _RAND_461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_462 = {1{`RANDOM}};
  _T_6887_399 = _RAND_462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_463 = {1{`RANDOM}};
  _T_6887_400 = _RAND_463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_464 = {1{`RANDOM}};
  _T_6887_401 = _RAND_464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_465 = {1{`RANDOM}};
  _T_6887_402 = _RAND_465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_466 = {1{`RANDOM}};
  _T_6887_403 = _RAND_466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_467 = {1{`RANDOM}};
  _T_6887_404 = _RAND_467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_468 = {1{`RANDOM}};
  _T_6887_405 = _RAND_468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_469 = {1{`RANDOM}};
  _T_6887_406 = _RAND_469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_470 = {1{`RANDOM}};
  _T_6887_407 = _RAND_470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_471 = {1{`RANDOM}};
  _T_6887_408 = _RAND_471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_472 = {1{`RANDOM}};
  _T_6887_409 = _RAND_472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_473 = {1{`RANDOM}};
  _T_6887_410 = _RAND_473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_474 = {1{`RANDOM}};
  _T_6887_411 = _RAND_474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_475 = {1{`RANDOM}};
  _T_6887_412 = _RAND_475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_476 = {1{`RANDOM}};
  _T_6887_413 = _RAND_476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_477 = {1{`RANDOM}};
  _T_6887_414 = _RAND_477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_478 = {1{`RANDOM}};
  _T_6887_415 = _RAND_478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_479 = {1{`RANDOM}};
  _T_6887_416 = _RAND_479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_480 = {1{`RANDOM}};
  _T_6887_417 = _RAND_480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_481 = {1{`RANDOM}};
  _T_6887_418 = _RAND_481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_482 = {1{`RANDOM}};
  _T_6887_419 = _RAND_482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_483 = {1{`RANDOM}};
  _T_6887_420 = _RAND_483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_484 = {1{`RANDOM}};
  _T_6887_421 = _RAND_484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_485 = {1{`RANDOM}};
  _T_6887_422 = _RAND_485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_486 = {1{`RANDOM}};
  _T_6887_423 = _RAND_486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_487 = {1{`RANDOM}};
  _T_6887_424 = _RAND_487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_488 = {1{`RANDOM}};
  _T_6887_425 = _RAND_488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_489 = {1{`RANDOM}};
  _T_6887_426 = _RAND_489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_490 = {1{`RANDOM}};
  _T_6887_427 = _RAND_490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_491 = {1{`RANDOM}};
  _T_6887_428 = _RAND_491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_492 = {1{`RANDOM}};
  _T_6887_429 = _RAND_492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_493 = {1{`RANDOM}};
  _T_6887_430 = _RAND_493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_494 = {1{`RANDOM}};
  _T_6887_431 = _RAND_494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_495 = {1{`RANDOM}};
  _T_6887_432 = _RAND_495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_496 = {1{`RANDOM}};
  _T_6887_433 = _RAND_496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_497 = {1{`RANDOM}};
  _T_6887_434 = _RAND_497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_498 = {1{`RANDOM}};
  _T_6887_435 = _RAND_498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_499 = {1{`RANDOM}};
  _T_6887_436 = _RAND_499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_500 = {1{`RANDOM}};
  _T_6887_437 = _RAND_500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_501 = {1{`RANDOM}};
  _T_6887_438 = _RAND_501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_502 = {1{`RANDOM}};
  _T_6887_439 = _RAND_502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_503 = {1{`RANDOM}};
  _T_6887_440 = _RAND_503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_504 = {1{`RANDOM}};
  _T_6887_441 = _RAND_504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_505 = {1{`RANDOM}};
  _T_6887_442 = _RAND_505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_506 = {1{`RANDOM}};
  _T_6887_443 = _RAND_506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_507 = {1{`RANDOM}};
  _T_6887_444 = _RAND_507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_508 = {1{`RANDOM}};
  _T_6887_445 = _RAND_508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_509 = {1{`RANDOM}};
  _T_6887_446 = _RAND_509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_510 = {1{`RANDOM}};
  _T_6887_447 = _RAND_510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_511 = {1{`RANDOM}};
  _T_6887_448 = _RAND_511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_512 = {1{`RANDOM}};
  _T_6887_449 = _RAND_512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_513 = {1{`RANDOM}};
  _T_6887_450 = _RAND_513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_514 = {1{`RANDOM}};
  _T_6887_451 = _RAND_514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_515 = {1{`RANDOM}};
  _T_6887_452 = _RAND_515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_516 = {1{`RANDOM}};
  _T_6887_453 = _RAND_516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_517 = {1{`RANDOM}};
  _T_6887_454 = _RAND_517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_518 = {1{`RANDOM}};
  _T_6887_455 = _RAND_518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_519 = {1{`RANDOM}};
  _T_6887_456 = _RAND_519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_520 = {1{`RANDOM}};
  _T_6887_457 = _RAND_520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_521 = {1{`RANDOM}};
  _T_6887_458 = _RAND_521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_522 = {1{`RANDOM}};
  _T_6887_459 = _RAND_522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_523 = {1{`RANDOM}};
  _T_6887_460 = _RAND_523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_524 = {1{`RANDOM}};
  _T_6887_461 = _RAND_524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_525 = {1{`RANDOM}};
  _T_6887_462 = _RAND_525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_526 = {1{`RANDOM}};
  _T_6887_463 = _RAND_526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_527 = {1{`RANDOM}};
  _T_6887_464 = _RAND_527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_528 = {1{`RANDOM}};
  _T_6887_465 = _RAND_528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_529 = {1{`RANDOM}};
  _T_6887_466 = _RAND_529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_530 = {1{`RANDOM}};
  _T_6887_467 = _RAND_530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_531 = {1{`RANDOM}};
  _T_6887_468 = _RAND_531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_532 = {1{`RANDOM}};
  _T_6887_469 = _RAND_532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_533 = {1{`RANDOM}};
  _T_6887_470 = _RAND_533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_534 = {1{`RANDOM}};
  _T_6887_471 = _RAND_534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_535 = {1{`RANDOM}};
  _T_6887_472 = _RAND_535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_536 = {1{`RANDOM}};
  _T_6887_473 = _RAND_536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_537 = {1{`RANDOM}};
  _T_6887_474 = _RAND_537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_538 = {1{`RANDOM}};
  _T_6887_475 = _RAND_538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_539 = {1{`RANDOM}};
  _T_6887_476 = _RAND_539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_540 = {1{`RANDOM}};
  _T_6887_477 = _RAND_540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_541 = {1{`RANDOM}};
  _T_6887_478 = _RAND_541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_542 = {1{`RANDOM}};
  _T_6887_479 = _RAND_542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_543 = {1{`RANDOM}};
  _T_6887_480 = _RAND_543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_544 = {1{`RANDOM}};
  _T_6887_481 = _RAND_544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_545 = {1{`RANDOM}};
  _T_6887_482 = _RAND_545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_546 = {1{`RANDOM}};
  _T_6887_483 = _RAND_546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_547 = {1{`RANDOM}};
  _T_6887_484 = _RAND_547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_548 = {1{`RANDOM}};
  _T_6887_485 = _RAND_548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_549 = {1{`RANDOM}};
  _T_6887_486 = _RAND_549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_550 = {1{`RANDOM}};
  _T_6887_487 = _RAND_550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_551 = {1{`RANDOM}};
  _T_6887_488 = _RAND_551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_552 = {1{`RANDOM}};
  _T_6887_489 = _RAND_552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_553 = {1{`RANDOM}};
  _T_6887_490 = _RAND_553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_554 = {1{`RANDOM}};
  _T_6887_491 = _RAND_554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_555 = {1{`RANDOM}};
  _T_6887_492 = _RAND_555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_556 = {1{`RANDOM}};
  _T_6887_493 = _RAND_556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_557 = {1{`RANDOM}};
  _T_6887_494 = _RAND_557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_558 = {1{`RANDOM}};
  _T_6887_495 = _RAND_558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_559 = {1{`RANDOM}};
  _T_6887_496 = _RAND_559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_560 = {1{`RANDOM}};
  _T_6887_497 = _RAND_560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_561 = {1{`RANDOM}};
  _T_6887_498 = _RAND_561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_562 = {1{`RANDOM}};
  _T_6887_499 = _RAND_562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_563 = {1{`RANDOM}};
  _T_6887_500 = _RAND_563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_564 = {1{`RANDOM}};
  _T_6887_501 = _RAND_564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_565 = {1{`RANDOM}};
  _T_6887_502 = _RAND_565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_566 = {1{`RANDOM}};
  _T_6887_503 = _RAND_566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_567 = {1{`RANDOM}};
  _T_6887_504 = _RAND_567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_568 = {1{`RANDOM}};
  _T_6887_505 = _RAND_568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_569 = {1{`RANDOM}};
  _T_6887_506 = _RAND_569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_570 = {1{`RANDOM}};
  _T_6887_507 = _RAND_570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_571 = {1{`RANDOM}};
  _T_6887_508 = _RAND_571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_572 = {1{`RANDOM}};
  _T_6887_509 = _RAND_572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_573 = {1{`RANDOM}};
  _T_6887_510 = _RAND_573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_574 = {1{`RANDOM}};
  _T_6887_511 = _RAND_574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_575 = {1{`RANDOM}};
  _T_6887_512 = _RAND_575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_576 = {1{`RANDOM}};
  _T_6887_513 = _RAND_576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_577 = {1{`RANDOM}};
  _T_6887_514 = _RAND_577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_578 = {1{`RANDOM}};
  _T_6887_515 = _RAND_578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_579 = {1{`RANDOM}};
  _T_6887_516 = _RAND_579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_580 = {1{`RANDOM}};
  _T_6887_517 = _RAND_580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_581 = {1{`RANDOM}};
  _T_6887_518 = _RAND_581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_582 = {1{`RANDOM}};
  _T_6887_519 = _RAND_582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_583 = {1{`RANDOM}};
  _T_6887_520 = _RAND_583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_584 = {1{`RANDOM}};
  _T_6887_521 = _RAND_584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_585 = {1{`RANDOM}};
  _T_6887_522 = _RAND_585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_586 = {1{`RANDOM}};
  _T_6887_523 = _RAND_586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_587 = {1{`RANDOM}};
  _T_6887_524 = _RAND_587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_588 = {1{`RANDOM}};
  _T_6887_525 = _RAND_588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_589 = {1{`RANDOM}};
  _T_6887_526 = _RAND_589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_590 = {1{`RANDOM}};
  _T_6887_527 = _RAND_590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_591 = {1{`RANDOM}};
  _T_6887_528 = _RAND_591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_592 = {1{`RANDOM}};
  _T_6887_529 = _RAND_592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_593 = {1{`RANDOM}};
  _T_6887_530 = _RAND_593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_594 = {1{`RANDOM}};
  _T_6887_531 = _RAND_594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_595 = {1{`RANDOM}};
  _T_6887_532 = _RAND_595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_596 = {1{`RANDOM}};
  _T_6887_533 = _RAND_596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_597 = {1{`RANDOM}};
  _T_6887_534 = _RAND_597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_598 = {1{`RANDOM}};
  _T_6887_535 = _RAND_598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_599 = {1{`RANDOM}};
  _T_6887_536 = _RAND_599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_600 = {1{`RANDOM}};
  _T_6887_537 = _RAND_600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_601 = {1{`RANDOM}};
  _T_6887_538 = _RAND_601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_602 = {1{`RANDOM}};
  _T_6887_539 = _RAND_602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_603 = {1{`RANDOM}};
  _T_6887_540 = _RAND_603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_604 = {1{`RANDOM}};
  _T_6887_541 = _RAND_604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_605 = {1{`RANDOM}};
  _T_6887_542 = _RAND_605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_606 = {1{`RANDOM}};
  _T_6887_543 = _RAND_606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_607 = {1{`RANDOM}};
  _T_6887_544 = _RAND_607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_608 = {1{`RANDOM}};
  _T_6887_545 = _RAND_608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_609 = {1{`RANDOM}};
  _T_6887_546 = _RAND_609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_610 = {1{`RANDOM}};
  _T_6887_547 = _RAND_610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_611 = {1{`RANDOM}};
  _T_6887_548 = _RAND_611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_612 = {1{`RANDOM}};
  _T_6887_549 = _RAND_612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_613 = {1{`RANDOM}};
  _T_6887_550 = _RAND_613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_614 = {1{`RANDOM}};
  _T_6887_551 = _RAND_614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_615 = {1{`RANDOM}};
  _T_6887_552 = _RAND_615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_616 = {1{`RANDOM}};
  _T_6887_553 = _RAND_616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_617 = {1{`RANDOM}};
  _T_6887_554 = _RAND_617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_618 = {1{`RANDOM}};
  _T_6887_555 = _RAND_618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_619 = {1{`RANDOM}};
  _T_6887_556 = _RAND_619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_620 = {1{`RANDOM}};
  _T_6887_557 = _RAND_620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_621 = {1{`RANDOM}};
  _T_6887_558 = _RAND_621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_622 = {1{`RANDOM}};
  _T_6887_559 = _RAND_622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_623 = {1{`RANDOM}};
  _T_6887_560 = _RAND_623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_624 = {1{`RANDOM}};
  _T_6887_561 = _RAND_624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_625 = {1{`RANDOM}};
  _T_6887_562 = _RAND_625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_626 = {1{`RANDOM}};
  _T_6887_563 = _RAND_626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_627 = {1{`RANDOM}};
  _T_6887_564 = _RAND_627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_628 = {1{`RANDOM}};
  _T_6887_565 = _RAND_628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_629 = {1{`RANDOM}};
  _T_6887_566 = _RAND_629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_630 = {1{`RANDOM}};
  _T_6887_567 = _RAND_630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_631 = {1{`RANDOM}};
  _T_6887_568 = _RAND_631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_632 = {1{`RANDOM}};
  _T_6887_569 = _RAND_632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_633 = {1{`RANDOM}};
  _T_6887_570 = _RAND_633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_634 = {1{`RANDOM}};
  _T_6887_571 = _RAND_634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_635 = {1{`RANDOM}};
  _T_6887_572 = _RAND_635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_636 = {1{`RANDOM}};
  _T_6887_573 = _RAND_636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_637 = {1{`RANDOM}};
  _T_6887_574 = _RAND_637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_638 = {1{`RANDOM}};
  _T_6887_575 = _RAND_638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_639 = {1{`RANDOM}};
  _T_6887_576 = _RAND_639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_640 = {1{`RANDOM}};
  _T_6887_577 = _RAND_640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_641 = {1{`RANDOM}};
  _T_6887_578 = _RAND_641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_642 = {1{`RANDOM}};
  _T_6887_579 = _RAND_642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_643 = {1{`RANDOM}};
  _T_6887_580 = _RAND_643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_644 = {1{`RANDOM}};
  _T_6887_581 = _RAND_644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_645 = {1{`RANDOM}};
  _T_6887_582 = _RAND_645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_646 = {1{`RANDOM}};
  _T_6887_583 = _RAND_646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_647 = {1{`RANDOM}};
  _T_6887_584 = _RAND_647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_648 = {1{`RANDOM}};
  _T_6887_585 = _RAND_648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_649 = {1{`RANDOM}};
  _T_6887_586 = _RAND_649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_650 = {1{`RANDOM}};
  _T_6887_587 = _RAND_650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_651 = {1{`RANDOM}};
  _T_6887_588 = _RAND_651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_652 = {1{`RANDOM}};
  _T_6887_589 = _RAND_652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_653 = {1{`RANDOM}};
  _T_6887_590 = _RAND_653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_654 = {1{`RANDOM}};
  _T_6887_591 = _RAND_654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_655 = {1{`RANDOM}};
  _T_6887_592 = _RAND_655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_656 = {1{`RANDOM}};
  _T_6887_593 = _RAND_656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_657 = {1{`RANDOM}};
  _T_6887_594 = _RAND_657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_658 = {1{`RANDOM}};
  _T_6887_595 = _RAND_658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_659 = {1{`RANDOM}};
  _T_6887_596 = _RAND_659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_660 = {1{`RANDOM}};
  _T_6887_597 = _RAND_660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_661 = {1{`RANDOM}};
  _T_6887_598 = _RAND_661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_662 = {1{`RANDOM}};
  _T_6887_599 = _RAND_662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_663 = {1{`RANDOM}};
  _T_6887_600 = _RAND_663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_664 = {1{`RANDOM}};
  _T_6887_601 = _RAND_664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_665 = {1{`RANDOM}};
  _T_6887_602 = _RAND_665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_666 = {1{`RANDOM}};
  _T_6887_603 = _RAND_666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_667 = {1{`RANDOM}};
  _T_6887_604 = _RAND_667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_668 = {1{`RANDOM}};
  _T_6887_605 = _RAND_668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_669 = {1{`RANDOM}};
  _T_6887_606 = _RAND_669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_670 = {1{`RANDOM}};
  _T_6887_607 = _RAND_670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_671 = {1{`RANDOM}};
  _T_6887_608 = _RAND_671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_672 = {1{`RANDOM}};
  _T_6887_609 = _RAND_672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_673 = {1{`RANDOM}};
  _T_6887_610 = _RAND_673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_674 = {1{`RANDOM}};
  _T_6887_611 = _RAND_674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_675 = {1{`RANDOM}};
  _T_6887_612 = _RAND_675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_676 = {1{`RANDOM}};
  _T_6887_613 = _RAND_676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_677 = {1{`RANDOM}};
  _T_6887_614 = _RAND_677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_678 = {1{`RANDOM}};
  _T_6887_615 = _RAND_678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_679 = {1{`RANDOM}};
  _T_6887_616 = _RAND_679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_680 = {1{`RANDOM}};
  _T_6887_617 = _RAND_680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_681 = {1{`RANDOM}};
  _T_6887_618 = _RAND_681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_682 = {1{`RANDOM}};
  _T_6887_619 = _RAND_682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_683 = {1{`RANDOM}};
  _T_6887_620 = _RAND_683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_684 = {1{`RANDOM}};
  _T_6887_621 = _RAND_684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_685 = {1{`RANDOM}};
  _T_6887_622 = _RAND_685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_686 = {1{`RANDOM}};
  _T_6887_623 = _RAND_686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_687 = {1{`RANDOM}};
  _T_6887_624 = _RAND_687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_688 = {1{`RANDOM}};
  _T_6887_625 = _RAND_688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_689 = {1{`RANDOM}};
  _T_6887_626 = _RAND_689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_690 = {1{`RANDOM}};
  _T_6887_627 = _RAND_690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_691 = {1{`RANDOM}};
  _T_6887_628 = _RAND_691[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_692 = {1{`RANDOM}};
  _T_6887_629 = _RAND_692[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_693 = {1{`RANDOM}};
  _T_6887_630 = _RAND_693[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_694 = {1{`RANDOM}};
  _T_6887_631 = _RAND_694[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_695 = {1{`RANDOM}};
  _T_6887_632 = _RAND_695[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_696 = {1{`RANDOM}};
  _T_6887_633 = _RAND_696[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_697 = {1{`RANDOM}};
  _T_6887_634 = _RAND_697[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_698 = {1{`RANDOM}};
  _T_6887_635 = _RAND_698[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_699 = {1{`RANDOM}};
  _T_6887_636 = _RAND_699[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_700 = {1{`RANDOM}};
  _T_6887_637 = _RAND_700[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_701 = {1{`RANDOM}};
  _T_6887_638 = _RAND_701[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_702 = {1{`RANDOM}};
  _T_6887_639 = _RAND_702[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_703 = {1{`RANDOM}};
  _T_6887_640 = _RAND_703[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_704 = {1{`RANDOM}};
  _T_6887_641 = _RAND_704[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_705 = {1{`RANDOM}};
  _T_6887_642 = _RAND_705[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_706 = {1{`RANDOM}};
  _T_6887_643 = _RAND_706[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_707 = {1{`RANDOM}};
  _T_6887_644 = _RAND_707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_708 = {1{`RANDOM}};
  _T_6887_645 = _RAND_708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_709 = {1{`RANDOM}};
  _T_6887_646 = _RAND_709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_710 = {1{`RANDOM}};
  _T_6887_647 = _RAND_710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_711 = {1{`RANDOM}};
  _T_6887_648 = _RAND_711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_712 = {1{`RANDOM}};
  _T_6887_649 = _RAND_712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_713 = {1{`RANDOM}};
  _T_6887_650 = _RAND_713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_714 = {1{`RANDOM}};
  _T_6887_651 = _RAND_714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_715 = {1{`RANDOM}};
  _T_6887_652 = _RAND_715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_716 = {1{`RANDOM}};
  _T_6887_653 = _RAND_716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_717 = {1{`RANDOM}};
  _T_6887_654 = _RAND_717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_718 = {1{`RANDOM}};
  _T_6887_655 = _RAND_718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_719 = {1{`RANDOM}};
  _T_6887_656 = _RAND_719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_720 = {1{`RANDOM}};
  _T_6887_657 = _RAND_720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_721 = {1{`RANDOM}};
  _T_6887_658 = _RAND_721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_722 = {1{`RANDOM}};
  _T_6887_659 = _RAND_722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_723 = {1{`RANDOM}};
  _T_6887_660 = _RAND_723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_724 = {1{`RANDOM}};
  _T_6887_661 = _RAND_724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_725 = {1{`RANDOM}};
  _T_6887_662 = _RAND_725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_726 = {1{`RANDOM}};
  _T_6887_663 = _RAND_726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_727 = {1{`RANDOM}};
  _T_6887_664 = _RAND_727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_728 = {1{`RANDOM}};
  _T_6887_665 = _RAND_728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_729 = {1{`RANDOM}};
  _T_6887_666 = _RAND_729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_730 = {1{`RANDOM}};
  _T_6887_667 = _RAND_730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_731 = {1{`RANDOM}};
  _T_6887_668 = _RAND_731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_732 = {1{`RANDOM}};
  _T_6887_669 = _RAND_732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_733 = {1{`RANDOM}};
  _T_6887_670 = _RAND_733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_734 = {1{`RANDOM}};
  _T_6887_671 = _RAND_734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_735 = {1{`RANDOM}};
  _T_6887_672 = _RAND_735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_736 = {1{`RANDOM}};
  _T_6887_673 = _RAND_736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_737 = {1{`RANDOM}};
  _T_6887_674 = _RAND_737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_738 = {1{`RANDOM}};
  _T_6887_675 = _RAND_738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_739 = {1{`RANDOM}};
  _T_6887_676 = _RAND_739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_740 = {1{`RANDOM}};
  _T_6887_677 = _RAND_740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_741 = {1{`RANDOM}};
  _T_6887_678 = _RAND_741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_742 = {1{`RANDOM}};
  _T_6887_679 = _RAND_742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_743 = {1{`RANDOM}};
  _T_6887_680 = _RAND_743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_744 = {1{`RANDOM}};
  _T_6887_681 = _RAND_744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_745 = {1{`RANDOM}};
  _T_6887_682 = _RAND_745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_746 = {1{`RANDOM}};
  _T_6887_683 = _RAND_746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_747 = {1{`RANDOM}};
  _T_6887_684 = _RAND_747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_748 = {1{`RANDOM}};
  _T_6887_685 = _RAND_748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_749 = {1{`RANDOM}};
  _T_6887_686 = _RAND_749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_750 = {1{`RANDOM}};
  _T_6887_687 = _RAND_750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_751 = {1{`RANDOM}};
  _T_6887_688 = _RAND_751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_752 = {1{`RANDOM}};
  _T_6887_689 = _RAND_752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_753 = {1{`RANDOM}};
  _T_6887_690 = _RAND_753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_754 = {1{`RANDOM}};
  _T_6887_691 = _RAND_754[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_755 = {1{`RANDOM}};
  _T_6887_692 = _RAND_755[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_756 = {1{`RANDOM}};
  _T_6887_693 = _RAND_756[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_757 = {1{`RANDOM}};
  _T_6887_694 = _RAND_757[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_758 = {1{`RANDOM}};
  _T_6887_695 = _RAND_758[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_759 = {1{`RANDOM}};
  _T_6887_696 = _RAND_759[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_760 = {1{`RANDOM}};
  _T_6887_697 = _RAND_760[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_761 = {1{`RANDOM}};
  _T_6887_698 = _RAND_761[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_762 = {1{`RANDOM}};
  _T_6887_699 = _RAND_762[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_763 = {1{`RANDOM}};
  _T_6887_700 = _RAND_763[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_764 = {1{`RANDOM}};
  _T_6887_701 = _RAND_764[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_765 = {1{`RANDOM}};
  _T_6887_702 = _RAND_765[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_766 = {1{`RANDOM}};
  _T_6887_703 = _RAND_766[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_767 = {1{`RANDOM}};
  _T_6887_704 = _RAND_767[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_768 = {1{`RANDOM}};
  _T_6887_705 = _RAND_768[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_769 = {1{`RANDOM}};
  _T_6887_706 = _RAND_769[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_770 = {1{`RANDOM}};
  _T_6887_707 = _RAND_770[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_771 = {1{`RANDOM}};
  _T_6887_708 = _RAND_771[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_772 = {1{`RANDOM}};
  _T_6887_709 = _RAND_772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_773 = {1{`RANDOM}};
  _T_6887_710 = _RAND_773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_774 = {1{`RANDOM}};
  _T_6887_711 = _RAND_774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_775 = {1{`RANDOM}};
  _T_6887_712 = _RAND_775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_776 = {1{`RANDOM}};
  _T_6887_713 = _RAND_776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_777 = {1{`RANDOM}};
  _T_6887_714 = _RAND_777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_778 = {1{`RANDOM}};
  _T_6887_715 = _RAND_778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_779 = {1{`RANDOM}};
  _T_6887_716 = _RAND_779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_780 = {1{`RANDOM}};
  _T_6887_717 = _RAND_780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_781 = {1{`RANDOM}};
  _T_6887_718 = _RAND_781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_782 = {1{`RANDOM}};
  _T_6887_719 = _RAND_782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_783 = {1{`RANDOM}};
  _T_6887_720 = _RAND_783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_784 = {1{`RANDOM}};
  _T_6887_721 = _RAND_784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_785 = {1{`RANDOM}};
  _T_6887_722 = _RAND_785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_786 = {1{`RANDOM}};
  _T_6887_723 = _RAND_786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_787 = {1{`RANDOM}};
  _T_6887_724 = _RAND_787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_788 = {1{`RANDOM}};
  _T_6887_725 = _RAND_788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_789 = {1{`RANDOM}};
  _T_6887_726 = _RAND_789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_790 = {1{`RANDOM}};
  _T_6887_727 = _RAND_790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_791 = {1{`RANDOM}};
  _T_6887_728 = _RAND_791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_792 = {1{`RANDOM}};
  _T_6887_729 = _RAND_792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_793 = {1{`RANDOM}};
  _T_6887_730 = _RAND_793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_794 = {1{`RANDOM}};
  _T_6887_731 = _RAND_794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_795 = {1{`RANDOM}};
  _T_6887_732 = _RAND_795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_796 = {1{`RANDOM}};
  _T_6887_733 = _RAND_796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_797 = {1{`RANDOM}};
  _T_6887_734 = _RAND_797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_798 = {1{`RANDOM}};
  _T_6887_735 = _RAND_798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_799 = {1{`RANDOM}};
  _T_6887_736 = _RAND_799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_800 = {1{`RANDOM}};
  _T_6887_737 = _RAND_800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_801 = {1{`RANDOM}};
  _T_6887_738 = _RAND_801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_802 = {1{`RANDOM}};
  _T_6887_739 = _RAND_802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_803 = {1{`RANDOM}};
  _T_6887_740 = _RAND_803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_804 = {1{`RANDOM}};
  _T_6887_741 = _RAND_804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_805 = {1{`RANDOM}};
  _T_6887_742 = _RAND_805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_806 = {1{`RANDOM}};
  _T_6887_743 = _RAND_806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_807 = {1{`RANDOM}};
  _T_6887_744 = _RAND_807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_808 = {1{`RANDOM}};
  _T_6887_745 = _RAND_808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_809 = {1{`RANDOM}};
  _T_6887_746 = _RAND_809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_810 = {1{`RANDOM}};
  _T_6887_747 = _RAND_810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_811 = {1{`RANDOM}};
  _T_6887_748 = _RAND_811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_812 = {1{`RANDOM}};
  _T_6887_749 = _RAND_812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_813 = {1{`RANDOM}};
  _T_6887_750 = _RAND_813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_814 = {1{`RANDOM}};
  _T_6887_751 = _RAND_814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_815 = {1{`RANDOM}};
  _T_6887_752 = _RAND_815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_816 = {1{`RANDOM}};
  _T_6887_753 = _RAND_816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_817 = {1{`RANDOM}};
  _T_6887_754 = _RAND_817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_818 = {1{`RANDOM}};
  _T_6887_755 = _RAND_818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_819 = {1{`RANDOM}};
  _T_6887_756 = _RAND_819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_820 = {1{`RANDOM}};
  _T_6887_757 = _RAND_820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_821 = {1{`RANDOM}};
  _T_6887_758 = _RAND_821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_822 = {1{`RANDOM}};
  _T_6887_759 = _RAND_822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_823 = {1{`RANDOM}};
  _T_6887_760 = _RAND_823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_824 = {1{`RANDOM}};
  _T_6887_761 = _RAND_824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_825 = {1{`RANDOM}};
  _T_6887_762 = _RAND_825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_826 = {1{`RANDOM}};
  _T_6887_763 = _RAND_826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_827 = {1{`RANDOM}};
  _T_6887_764 = _RAND_827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_828 = {1{`RANDOM}};
  _T_6887_765 = _RAND_828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_829 = {1{`RANDOM}};
  _T_6887_766 = _RAND_829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_830 = {1{`RANDOM}};
  _T_6887_767 = _RAND_830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_831 = {1{`RANDOM}};
  _T_6887_768 = _RAND_831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_832 = {1{`RANDOM}};
  _T_6887_769 = _RAND_832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_833 = {1{`RANDOM}};
  _T_6887_770 = _RAND_833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_834 = {1{`RANDOM}};
  _T_6887_771 = _RAND_834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_835 = {1{`RANDOM}};
  _T_6887_772 = _RAND_835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_836 = {1{`RANDOM}};
  _T_6887_773 = _RAND_836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_837 = {1{`RANDOM}};
  _T_6887_774 = _RAND_837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_838 = {1{`RANDOM}};
  _T_6887_775 = _RAND_838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_839 = {1{`RANDOM}};
  _T_6887_776 = _RAND_839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_840 = {1{`RANDOM}};
  _T_6887_777 = _RAND_840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_841 = {1{`RANDOM}};
  _T_6887_778 = _RAND_841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_842 = {1{`RANDOM}};
  _T_6887_779 = _RAND_842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_843 = {1{`RANDOM}};
  _T_6887_780 = _RAND_843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_844 = {1{`RANDOM}};
  _T_6887_781 = _RAND_844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_845 = {1{`RANDOM}};
  _T_6887_782 = _RAND_845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_846 = {1{`RANDOM}};
  _T_6887_783 = _RAND_846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_847 = {1{`RANDOM}};
  _T_6887_784 = _RAND_847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_848 = {1{`RANDOM}};
  _T_6887_785 = _RAND_848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_849 = {1{`RANDOM}};
  _T_6887_786 = _RAND_849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_850 = {1{`RANDOM}};
  _T_6887_787 = _RAND_850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_851 = {1{`RANDOM}};
  _T_6887_788 = _RAND_851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_852 = {1{`RANDOM}};
  _T_6887_789 = _RAND_852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_853 = {1{`RANDOM}};
  _T_6887_790 = _RAND_853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_854 = {1{`RANDOM}};
  _T_6887_791 = _RAND_854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_855 = {1{`RANDOM}};
  _T_6887_792 = _RAND_855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_856 = {1{`RANDOM}};
  _T_6887_793 = _RAND_856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_857 = {1{`RANDOM}};
  _T_6887_794 = _RAND_857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_858 = {1{`RANDOM}};
  _T_6887_795 = _RAND_858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_859 = {1{`RANDOM}};
  _T_6887_796 = _RAND_859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_860 = {1{`RANDOM}};
  _T_6887_797 = _RAND_860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_861 = {1{`RANDOM}};
  _T_6887_798 = _RAND_861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_862 = {1{`RANDOM}};
  _T_6887_799 = _RAND_862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_863 = {1{`RANDOM}};
  _T_6887_800 = _RAND_863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_864 = {1{`RANDOM}};
  _T_6887_801 = _RAND_864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_865 = {1{`RANDOM}};
  _T_6887_802 = _RAND_865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_866 = {1{`RANDOM}};
  _T_6887_803 = _RAND_866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_867 = {1{`RANDOM}};
  _T_6887_804 = _RAND_867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_868 = {1{`RANDOM}};
  _T_6887_805 = _RAND_868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_869 = {1{`RANDOM}};
  _T_6887_806 = _RAND_869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_870 = {1{`RANDOM}};
  _T_6887_807 = _RAND_870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_871 = {1{`RANDOM}};
  _T_6887_808 = _RAND_871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_872 = {1{`RANDOM}};
  _T_6887_809 = _RAND_872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_873 = {1{`RANDOM}};
  _T_6887_810 = _RAND_873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_874 = {1{`RANDOM}};
  _T_6887_811 = _RAND_874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_875 = {1{`RANDOM}};
  _T_6887_812 = _RAND_875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_876 = {1{`RANDOM}};
  _T_6887_813 = _RAND_876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_877 = {1{`RANDOM}};
  _T_6887_814 = _RAND_877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_878 = {1{`RANDOM}};
  _T_6887_815 = _RAND_878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_879 = {1{`RANDOM}};
  _T_6887_816 = _RAND_879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_880 = {1{`RANDOM}};
  _T_6887_817 = _RAND_880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_881 = {1{`RANDOM}};
  _T_6887_818 = _RAND_881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_882 = {1{`RANDOM}};
  _T_6887_819 = _RAND_882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_883 = {1{`RANDOM}};
  _T_6887_820 = _RAND_883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_884 = {1{`RANDOM}};
  _T_6887_821 = _RAND_884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_885 = {1{`RANDOM}};
  _T_6887_822 = _RAND_885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_886 = {1{`RANDOM}};
  _T_6887_823 = _RAND_886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_887 = {1{`RANDOM}};
  _T_6887_824 = _RAND_887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_888 = {1{`RANDOM}};
  _T_6887_825 = _RAND_888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_889 = {1{`RANDOM}};
  _T_6887_826 = _RAND_889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_890 = {1{`RANDOM}};
  _T_6887_827 = _RAND_890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_891 = {1{`RANDOM}};
  _T_6887_828 = _RAND_891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_892 = {1{`RANDOM}};
  _T_6887_829 = _RAND_892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_893 = {1{`RANDOM}};
  _T_6887_830 = _RAND_893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_894 = {1{`RANDOM}};
  _T_6887_831 = _RAND_894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_895 = {1{`RANDOM}};
  _T_6887_832 = _RAND_895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_896 = {1{`RANDOM}};
  _T_6887_833 = _RAND_896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_897 = {1{`RANDOM}};
  _T_6887_834 = _RAND_897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_898 = {1{`RANDOM}};
  _T_6887_835 = _RAND_898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_899 = {1{`RANDOM}};
  _T_6887_836 = _RAND_899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_900 = {1{`RANDOM}};
  _T_6887_837 = _RAND_900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_901 = {1{`RANDOM}};
  _T_6887_838 = _RAND_901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_902 = {1{`RANDOM}};
  _T_6887_839 = _RAND_902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_903 = {1{`RANDOM}};
  _T_6887_840 = _RAND_903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_904 = {1{`RANDOM}};
  _T_6887_841 = _RAND_904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_905 = {1{`RANDOM}};
  _T_6887_842 = _RAND_905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_906 = {1{`RANDOM}};
  _T_6887_843 = _RAND_906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_907 = {1{`RANDOM}};
  _T_6887_844 = _RAND_907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_908 = {1{`RANDOM}};
  _T_6887_845 = _RAND_908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_909 = {1{`RANDOM}};
  _T_6887_846 = _RAND_909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_910 = {1{`RANDOM}};
  _T_6887_847 = _RAND_910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_911 = {1{`RANDOM}};
  _T_6887_848 = _RAND_911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_912 = {1{`RANDOM}};
  _T_6887_849 = _RAND_912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_913 = {1{`RANDOM}};
  _T_6887_850 = _RAND_913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_914 = {1{`RANDOM}};
  _T_6887_851 = _RAND_914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_915 = {1{`RANDOM}};
  _T_6887_852 = _RAND_915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_916 = {1{`RANDOM}};
  _T_6887_853 = _RAND_916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_917 = {1{`RANDOM}};
  _T_6887_854 = _RAND_917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_918 = {1{`RANDOM}};
  _T_6887_855 = _RAND_918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_919 = {1{`RANDOM}};
  _T_6887_856 = _RAND_919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_920 = {1{`RANDOM}};
  _T_6887_857 = _RAND_920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_921 = {1{`RANDOM}};
  _T_6887_858 = _RAND_921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_922 = {1{`RANDOM}};
  _T_6887_859 = _RAND_922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_923 = {1{`RANDOM}};
  _T_6887_860 = _RAND_923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_924 = {1{`RANDOM}};
  _T_6887_861 = _RAND_924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_925 = {1{`RANDOM}};
  _T_6887_862 = _RAND_925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_926 = {1{`RANDOM}};
  _T_6887_863 = _RAND_926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_927 = {1{`RANDOM}};
  _T_6887_864 = _RAND_927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_928 = {1{`RANDOM}};
  _T_6887_865 = _RAND_928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_929 = {1{`RANDOM}};
  _T_6887_866 = _RAND_929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_930 = {1{`RANDOM}};
  _T_6887_867 = _RAND_930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_931 = {1{`RANDOM}};
  _T_6887_868 = _RAND_931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_932 = {1{`RANDOM}};
  _T_6887_869 = _RAND_932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_933 = {1{`RANDOM}};
  _T_6887_870 = _RAND_933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_934 = {1{`RANDOM}};
  _T_6887_871 = _RAND_934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_935 = {1{`RANDOM}};
  _T_6887_872 = _RAND_935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_936 = {1{`RANDOM}};
  _T_6887_873 = _RAND_936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_937 = {1{`RANDOM}};
  _T_6887_874 = _RAND_937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_938 = {1{`RANDOM}};
  _T_6887_875 = _RAND_938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_939 = {1{`RANDOM}};
  _T_6887_876 = _RAND_939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_940 = {1{`RANDOM}};
  _T_6887_877 = _RAND_940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_941 = {1{`RANDOM}};
  _T_6887_878 = _RAND_941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_942 = {1{`RANDOM}};
  _T_6887_879 = _RAND_942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_943 = {1{`RANDOM}};
  _T_6887_880 = _RAND_943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_944 = {1{`RANDOM}};
  _T_6887_881 = _RAND_944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_945 = {1{`RANDOM}};
  _T_6887_882 = _RAND_945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_946 = {1{`RANDOM}};
  _T_6887_883 = _RAND_946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_947 = {1{`RANDOM}};
  _T_6887_884 = _RAND_947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_948 = {1{`RANDOM}};
  _T_6887_885 = _RAND_948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_949 = {1{`RANDOM}};
  _T_6887_886 = _RAND_949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_950 = {1{`RANDOM}};
  _T_6887_887 = _RAND_950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_951 = {1{`RANDOM}};
  _T_6887_888 = _RAND_951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_952 = {1{`RANDOM}};
  _T_6887_889 = _RAND_952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_953 = {1{`RANDOM}};
  _T_6887_890 = _RAND_953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_954 = {1{`RANDOM}};
  _T_6887_891 = _RAND_954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_955 = {1{`RANDOM}};
  _T_6887_892 = _RAND_955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_956 = {1{`RANDOM}};
  _T_6887_893 = _RAND_956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_957 = {1{`RANDOM}};
  _T_6887_894 = _RAND_957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_958 = {1{`RANDOM}};
  _T_6887_895 = _RAND_958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_959 = {1{`RANDOM}};
  _T_6887_896 = _RAND_959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_960 = {1{`RANDOM}};
  _T_6887_897 = _RAND_960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_961 = {1{`RANDOM}};
  _T_6887_898 = _RAND_961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_962 = {1{`RANDOM}};
  _T_6887_899 = _RAND_962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_963 = {1{`RANDOM}};
  _T_6887_900 = _RAND_963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_964 = {1{`RANDOM}};
  _T_6887_901 = _RAND_964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_965 = {1{`RANDOM}};
  _T_6887_902 = _RAND_965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_966 = {1{`RANDOM}};
  _T_6887_903 = _RAND_966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_967 = {1{`RANDOM}};
  _T_6887_904 = _RAND_967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_968 = {1{`RANDOM}};
  _T_6887_905 = _RAND_968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_969 = {1{`RANDOM}};
  _T_6887_906 = _RAND_969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_970 = {1{`RANDOM}};
  _T_6887_907 = _RAND_970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_971 = {1{`RANDOM}};
  _T_6887_908 = _RAND_971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_972 = {1{`RANDOM}};
  _T_6887_909 = _RAND_972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_973 = {1{`RANDOM}};
  _T_6887_910 = _RAND_973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_974 = {1{`RANDOM}};
  _T_6887_911 = _RAND_974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_975 = {1{`RANDOM}};
  _T_6887_912 = _RAND_975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_976 = {1{`RANDOM}};
  _T_6887_913 = _RAND_976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_977 = {1{`RANDOM}};
  _T_6887_914 = _RAND_977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_978 = {1{`RANDOM}};
  _T_6887_915 = _RAND_978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_979 = {1{`RANDOM}};
  _T_6887_916 = _RAND_979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_980 = {1{`RANDOM}};
  _T_6887_917 = _RAND_980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_981 = {1{`RANDOM}};
  _T_6887_918 = _RAND_981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_982 = {1{`RANDOM}};
  _T_6887_919 = _RAND_982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_983 = {1{`RANDOM}};
  _T_6887_920 = _RAND_983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_984 = {1{`RANDOM}};
  _T_6887_921 = _RAND_984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_985 = {1{`RANDOM}};
  _T_6887_922 = _RAND_985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_986 = {1{`RANDOM}};
  _T_6887_923 = _RAND_986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_987 = {1{`RANDOM}};
  _T_6887_924 = _RAND_987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_988 = {1{`RANDOM}};
  _T_6887_925 = _RAND_988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_989 = {1{`RANDOM}};
  _T_6887_926 = _RAND_989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_990 = {1{`RANDOM}};
  _T_6887_927 = _RAND_990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_991 = {1{`RANDOM}};
  _T_6887_928 = _RAND_991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_992 = {1{`RANDOM}};
  _T_6887_929 = _RAND_992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_993 = {1{`RANDOM}};
  _T_6887_930 = _RAND_993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_994 = {1{`RANDOM}};
  _T_6887_931 = _RAND_994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_995 = {1{`RANDOM}};
  _T_6887_932 = _RAND_995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_996 = {1{`RANDOM}};
  _T_6887_933 = _RAND_996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_997 = {1{`RANDOM}};
  _T_6887_934 = _RAND_997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_998 = {1{`RANDOM}};
  _T_6887_935 = _RAND_998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_999 = {1{`RANDOM}};
  _T_6887_936 = _RAND_999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1000 = {1{`RANDOM}};
  _T_6887_937 = _RAND_1000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1001 = {1{`RANDOM}};
  _T_6887_938 = _RAND_1001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1002 = {1{`RANDOM}};
  _T_6887_939 = _RAND_1002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1003 = {1{`RANDOM}};
  _T_6887_940 = _RAND_1003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1004 = {1{`RANDOM}};
  _T_6887_941 = _RAND_1004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1005 = {1{`RANDOM}};
  _T_6887_942 = _RAND_1005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1006 = {1{`RANDOM}};
  _T_6887_943 = _RAND_1006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1007 = {1{`RANDOM}};
  _T_6887_944 = _RAND_1007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1008 = {1{`RANDOM}};
  _T_6887_945 = _RAND_1008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1009 = {1{`RANDOM}};
  _T_6887_946 = _RAND_1009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1010 = {1{`RANDOM}};
  _T_6887_947 = _RAND_1010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1011 = {1{`RANDOM}};
  _T_6887_948 = _RAND_1011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1012 = {1{`RANDOM}};
  _T_6887_949 = _RAND_1012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1013 = {1{`RANDOM}};
  _T_6887_950 = _RAND_1013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1014 = {1{`RANDOM}};
  _T_6887_951 = _RAND_1014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1015 = {1{`RANDOM}};
  _T_6887_952 = _RAND_1015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1016 = {1{`RANDOM}};
  _T_6887_953 = _RAND_1016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1017 = {1{`RANDOM}};
  _T_6887_954 = _RAND_1017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1018 = {1{`RANDOM}};
  _T_6887_955 = _RAND_1018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1019 = {1{`RANDOM}};
  _T_6887_956 = _RAND_1019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1020 = {1{`RANDOM}};
  _T_6887_957 = _RAND_1020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1021 = {1{`RANDOM}};
  _T_6887_958 = _RAND_1021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1022 = {1{`RANDOM}};
  _T_6887_959 = _RAND_1022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1023 = {1{`RANDOM}};
  _T_6887_960 = _RAND_1023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1024 = {1{`RANDOM}};
  _T_6887_961 = _RAND_1024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1025 = {1{`RANDOM}};
  _T_6887_962 = _RAND_1025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1026 = {1{`RANDOM}};
  _T_6887_963 = _RAND_1026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1027 = {1{`RANDOM}};
  _T_6887_964 = _RAND_1027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1028 = {1{`RANDOM}};
  _T_6887_965 = _RAND_1028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1029 = {1{`RANDOM}};
  _T_6887_966 = _RAND_1029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1030 = {1{`RANDOM}};
  _T_6887_967 = _RAND_1030[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1031 = {1{`RANDOM}};
  _T_6887_968 = _RAND_1031[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1032 = {1{`RANDOM}};
  _T_6887_969 = _RAND_1032[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1033 = {1{`RANDOM}};
  _T_6887_970 = _RAND_1033[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1034 = {1{`RANDOM}};
  _T_6887_971 = _RAND_1034[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1035 = {1{`RANDOM}};
  _T_6887_972 = _RAND_1035[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1036 = {1{`RANDOM}};
  _T_6887_973 = _RAND_1036[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1037 = {1{`RANDOM}};
  _T_6887_974 = _RAND_1037[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1038 = {1{`RANDOM}};
  _T_6887_975 = _RAND_1038[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1039 = {1{`RANDOM}};
  _T_6887_976 = _RAND_1039[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1040 = {1{`RANDOM}};
  _T_6887_977 = _RAND_1040[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1041 = {1{`RANDOM}};
  _T_6887_978 = _RAND_1041[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1042 = {1{`RANDOM}};
  _T_6887_979 = _RAND_1042[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1043 = {1{`RANDOM}};
  _T_6887_980 = _RAND_1043[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1044 = {1{`RANDOM}};
  _T_6887_981 = _RAND_1044[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1045 = {1{`RANDOM}};
  _T_6887_982 = _RAND_1045[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1046 = {1{`RANDOM}};
  _T_6887_983 = _RAND_1046[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1047 = {1{`RANDOM}};
  _T_6887_984 = _RAND_1047[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1048 = {1{`RANDOM}};
  _T_6887_985 = _RAND_1048[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1049 = {1{`RANDOM}};
  _T_6887_986 = _RAND_1049[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1050 = {1{`RANDOM}};
  _T_6887_987 = _RAND_1050[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1051 = {1{`RANDOM}};
  _T_6887_988 = _RAND_1051[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1052 = {1{`RANDOM}};
  _T_6887_989 = _RAND_1052[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1053 = {1{`RANDOM}};
  _T_6887_990 = _RAND_1053[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1054 = {1{`RANDOM}};
  _T_6887_991 = _RAND_1054[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1055 = {1{`RANDOM}};
  _T_6887_992 = _RAND_1055[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1056 = {1{`RANDOM}};
  _T_6887_993 = _RAND_1056[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1057 = {1{`RANDOM}};
  _T_6887_994 = _RAND_1057[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1058 = {1{`RANDOM}};
  _T_6887_995 = _RAND_1058[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1059 = {1{`RANDOM}};
  _T_6887_996 = _RAND_1059[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1060 = {1{`RANDOM}};
  _T_6887_997 = _RAND_1060[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1061 = {1{`RANDOM}};
  _T_6887_998 = _RAND_1061[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1062 = {1{`RANDOM}};
  _T_6887_999 = _RAND_1062[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1063 = {1{`RANDOM}};
  _T_6887_1000 = _RAND_1063[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1064 = {1{`RANDOM}};
  _T_6887_1001 = _RAND_1064[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1065 = {1{`RANDOM}};
  _T_6887_1002 = _RAND_1065[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1066 = {1{`RANDOM}};
  _T_6887_1003 = _RAND_1066[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1067 = {1{`RANDOM}};
  _T_6887_1004 = _RAND_1067[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1068 = {1{`RANDOM}};
  _T_6887_1005 = _RAND_1068[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1069 = {1{`RANDOM}};
  _T_6887_1006 = _RAND_1069[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1070 = {1{`RANDOM}};
  _T_6887_1007 = _RAND_1070[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1071 = {1{`RANDOM}};
  _T_6887_1008 = _RAND_1071[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1072 = {1{`RANDOM}};
  _T_6887_1009 = _RAND_1072[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1073 = {1{`RANDOM}};
  _T_6887_1010 = _RAND_1073[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1074 = {1{`RANDOM}};
  _T_6887_1011 = _RAND_1074[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1075 = {1{`RANDOM}};
  _T_6887_1012 = _RAND_1075[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1076 = {1{`RANDOM}};
  _T_6887_1013 = _RAND_1076[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1077 = {1{`RANDOM}};
  _T_6887_1014 = _RAND_1077[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1078 = {1{`RANDOM}};
  _T_6887_1015 = _RAND_1078[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1079 = {1{`RANDOM}};
  _T_6887_1016 = _RAND_1079[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1080 = {1{`RANDOM}};
  _T_6887_1017 = _RAND_1080[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1081 = {1{`RANDOM}};
  _T_6887_1018 = _RAND_1081[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1082 = {1{`RANDOM}};
  _T_6887_1019 = _RAND_1082[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1083 = {1{`RANDOM}};
  _T_6887_1020 = _RAND_1083[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1084 = {1{`RANDOM}};
  _T_6887_1021 = _RAND_1084[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1085 = {1{`RANDOM}};
  _T_6887_1022 = _RAND_1085[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1086 = {1{`RANDOM}};
  _T_6887_1023 = _RAND_1086[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1087 = {1{`RANDOM}};
  _T_6887_1024 = _RAND_1087[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1088 = {1{`RANDOM}};
  _T_6887_1025 = _RAND_1088[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1089 = {1{`RANDOM}};
  _T_6887_1026 = _RAND_1089[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1090 = {1{`RANDOM}};
  _T_6887_1027 = _RAND_1090[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1091 = {1{`RANDOM}};
  _T_6887_1028 = _RAND_1091[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1092 = {1{`RANDOM}};
  _T_6887_1029 = _RAND_1092[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1093 = {1{`RANDOM}};
  _T_6887_1030 = _RAND_1093[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1094 = {1{`RANDOM}};
  _T_6887_1031 = _RAND_1094[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1095 = {1{`RANDOM}};
  _T_6887_1032 = _RAND_1095[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1096 = {1{`RANDOM}};
  _T_6887_1033 = _RAND_1096[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1097 = {1{`RANDOM}};
  _T_6887_1034 = _RAND_1097[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1098 = {1{`RANDOM}};
  _T_6887_1035 = _RAND_1098[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1099 = {1{`RANDOM}};
  _T_6887_1036 = _RAND_1099[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1100 = {1{`RANDOM}};
  _T_6887_1037 = _RAND_1100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1101 = {1{`RANDOM}};
  _T_6887_1038 = _RAND_1101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1102 = {1{`RANDOM}};
  _T_6887_1039 = _RAND_1102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1103 = {1{`RANDOM}};
  _T_6887_1040 = _RAND_1103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1104 = {1{`RANDOM}};
  _T_6887_1041 = _RAND_1104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1105 = {1{`RANDOM}};
  _T_6887_1042 = _RAND_1105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1106 = {1{`RANDOM}};
  _T_6887_1043 = _RAND_1106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1107 = {1{`RANDOM}};
  _T_6887_1044 = _RAND_1107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1108 = {1{`RANDOM}};
  _T_6887_1045 = _RAND_1108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1109 = {1{`RANDOM}};
  _T_6887_1046 = _RAND_1109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1110 = {1{`RANDOM}};
  _T_6887_1047 = _RAND_1110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1111 = {1{`RANDOM}};
  _T_6887_1048 = _RAND_1111[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1112 = {1{`RANDOM}};
  _T_6887_1049 = _RAND_1112[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1113 = {1{`RANDOM}};
  _T_6887_1050 = _RAND_1113[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1114 = {1{`RANDOM}};
  _T_6887_1051 = _RAND_1114[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1115 = {1{`RANDOM}};
  _T_6887_1052 = _RAND_1115[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1116 = {1{`RANDOM}};
  _T_6887_1053 = _RAND_1116[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1117 = {1{`RANDOM}};
  _T_6887_1054 = _RAND_1117[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1118 = {1{`RANDOM}};
  _T_6887_1055 = _RAND_1118[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1119 = {1{`RANDOM}};
  _T_6887_1056 = _RAND_1119[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1120 = {1{`RANDOM}};
  _T_6887_1057 = _RAND_1120[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1121 = {1{`RANDOM}};
  _T_6887_1058 = _RAND_1121[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1122 = {1{`RANDOM}};
  _T_6887_1059 = _RAND_1122[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1123 = {1{`RANDOM}};
  _T_6887_1060 = _RAND_1123[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1124 = {1{`RANDOM}};
  _T_6887_1061 = _RAND_1124[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1125 = {1{`RANDOM}};
  _T_6887_1062 = _RAND_1125[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1126 = {1{`RANDOM}};
  _T_6887_1063 = _RAND_1126[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1127 = {1{`RANDOM}};
  _T_6887_1064 = _RAND_1127[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1128 = {1{`RANDOM}};
  _T_6887_1065 = _RAND_1128[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1129 = {1{`RANDOM}};
  _T_6887_1066 = _RAND_1129[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1130 = {1{`RANDOM}};
  _T_6887_1067 = _RAND_1130[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1131 = {1{`RANDOM}};
  _T_6887_1068 = _RAND_1131[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1132 = {1{`RANDOM}};
  _T_6887_1069 = _RAND_1132[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1133 = {1{`RANDOM}};
  _T_6887_1070 = _RAND_1133[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1134 = {1{`RANDOM}};
  _T_6887_1071 = _RAND_1134[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1135 = {1{`RANDOM}};
  _T_6887_1072 = _RAND_1135[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1136 = {1{`RANDOM}};
  _T_6887_1073 = _RAND_1136[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1137 = {1{`RANDOM}};
  _T_6887_1074 = _RAND_1137[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1138 = {1{`RANDOM}};
  _T_6887_1075 = _RAND_1138[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1139 = {1{`RANDOM}};
  _T_6887_1076 = _RAND_1139[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1140 = {1{`RANDOM}};
  _T_6887_1077 = _RAND_1140[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1141 = {1{`RANDOM}};
  _T_6887_1078 = _RAND_1141[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1142 = {1{`RANDOM}};
  _T_6887_1079 = _RAND_1142[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1143 = {1{`RANDOM}};
  _T_6887_1080 = _RAND_1143[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1144 = {1{`RANDOM}};
  _T_6887_1081 = _RAND_1144[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1145 = {1{`RANDOM}};
  _T_6887_1082 = _RAND_1145[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1146 = {1{`RANDOM}};
  _T_6887_1083 = _RAND_1146[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1147 = {1{`RANDOM}};
  _T_6887_1084 = _RAND_1147[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1148 = {1{`RANDOM}};
  _T_6887_1085 = _RAND_1148[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1149 = {1{`RANDOM}};
  _T_6887_1086 = _RAND_1149[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1150 = {1{`RANDOM}};
  _T_6887_1087 = _RAND_1150[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1151 = {1{`RANDOM}};
  _T_6887_1088 = _RAND_1151[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1152 = {1{`RANDOM}};
  _T_6887_1089 = _RAND_1152[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1153 = {1{`RANDOM}};
  _T_6887_1090 = _RAND_1153[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1154 = {1{`RANDOM}};
  _T_6887_1091 = _RAND_1154[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1155 = {1{`RANDOM}};
  _T_6887_1092 = _RAND_1155[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1156 = {1{`RANDOM}};
  _T_6887_1093 = _RAND_1156[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1157 = {1{`RANDOM}};
  _T_6887_1094 = _RAND_1157[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1158 = {1{`RANDOM}};
  _T_6887_1095 = _RAND_1158[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1159 = {1{`RANDOM}};
  _T_6887_1096 = _RAND_1159[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1160 = {1{`RANDOM}};
  _T_6887_1097 = _RAND_1160[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1161 = {1{`RANDOM}};
  _T_6887_1098 = _RAND_1161[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1162 = {1{`RANDOM}};
  _T_6887_1099 = _RAND_1162[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1163 = {1{`RANDOM}};
  _T_6887_1100 = _RAND_1163[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1164 = {1{`RANDOM}};
  _T_6887_1101 = _RAND_1164[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1165 = {1{`RANDOM}};
  _T_6887_1102 = _RAND_1165[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1166 = {1{`RANDOM}};
  _T_6887_1103 = _RAND_1166[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1167 = {1{`RANDOM}};
  _T_6887_1104 = _RAND_1167[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1168 = {1{`RANDOM}};
  _T_6887_1105 = _RAND_1168[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1169 = {1{`RANDOM}};
  _T_6887_1106 = _RAND_1169[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1170 = {1{`RANDOM}};
  _T_6887_1107 = _RAND_1170[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1171 = {1{`RANDOM}};
  _T_6887_1108 = _RAND_1171[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1172 = {1{`RANDOM}};
  _T_6887_1109 = _RAND_1172[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1173 = {1{`RANDOM}};
  _T_6887_1110 = _RAND_1173[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1174 = {1{`RANDOM}};
  _T_6887_1111 = _RAND_1174[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1175 = {1{`RANDOM}};
  _T_6887_1112 = _RAND_1175[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1176 = {1{`RANDOM}};
  _T_6887_1113 = _RAND_1176[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1177 = {1{`RANDOM}};
  _T_6887_1114 = _RAND_1177[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1178 = {1{`RANDOM}};
  _T_6887_1115 = _RAND_1178[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1179 = {1{`RANDOM}};
  _T_6887_1116 = _RAND_1179[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1180 = {1{`RANDOM}};
  _T_6887_1117 = _RAND_1180[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1181 = {1{`RANDOM}};
  _T_6887_1118 = _RAND_1181[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1182 = {1{`RANDOM}};
  _T_6887_1119 = _RAND_1182[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1183 = {1{`RANDOM}};
  _T_6887_1120 = _RAND_1183[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1184 = {1{`RANDOM}};
  _T_6887_1121 = _RAND_1184[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1185 = {1{`RANDOM}};
  _T_6887_1122 = _RAND_1185[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1186 = {1{`RANDOM}};
  _T_6887_1123 = _RAND_1186[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1187 = {1{`RANDOM}};
  _T_6887_1124 = _RAND_1187[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1188 = {1{`RANDOM}};
  _T_6887_1125 = _RAND_1188[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1189 = {1{`RANDOM}};
  _T_6887_1126 = _RAND_1189[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1190 = {1{`RANDOM}};
  _T_6887_1127 = _RAND_1190[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1191 = {1{`RANDOM}};
  _T_6887_1128 = _RAND_1191[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1192 = {1{`RANDOM}};
  _T_6887_1129 = _RAND_1192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1193 = {1{`RANDOM}};
  _T_6887_1130 = _RAND_1193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1194 = {1{`RANDOM}};
  _T_6887_1131 = _RAND_1194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1195 = {1{`RANDOM}};
  _T_6887_1132 = _RAND_1195[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1196 = {1{`RANDOM}};
  _T_6887_1133 = _RAND_1196[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1197 = {1{`RANDOM}};
  _T_6887_1134 = _RAND_1197[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1198 = {1{`RANDOM}};
  _T_6887_1135 = _RAND_1198[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1199 = {1{`RANDOM}};
  _T_6887_1136 = _RAND_1199[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1200 = {1{`RANDOM}};
  _T_6887_1137 = _RAND_1200[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1201 = {1{`RANDOM}};
  _T_6887_1138 = _RAND_1201[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1202 = {1{`RANDOM}};
  _T_6887_1139 = _RAND_1202[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1203 = {1{`RANDOM}};
  _T_6887_1140 = _RAND_1203[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1204 = {1{`RANDOM}};
  _T_6887_1141 = _RAND_1204[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1205 = {1{`RANDOM}};
  _T_6887_1142 = _RAND_1205[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1206 = {1{`RANDOM}};
  _T_6887_1143 = _RAND_1206[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1207 = {1{`RANDOM}};
  _T_6887_1144 = _RAND_1207[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1208 = {1{`RANDOM}};
  _T_6887_1145 = _RAND_1208[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1209 = {1{`RANDOM}};
  _T_6887_1146 = _RAND_1209[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1210 = {1{`RANDOM}};
  _T_6887_1147 = _RAND_1210[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1211 = {1{`RANDOM}};
  _T_6887_1148 = _RAND_1211[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1212 = {1{`RANDOM}};
  _T_6887_1149 = _RAND_1212[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1213 = {1{`RANDOM}};
  _T_6887_1150 = _RAND_1213[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1214 = {1{`RANDOM}};
  _T_6887_1151 = _RAND_1214[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1215 = {1{`RANDOM}};
  _T_6887_1152 = _RAND_1215[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1216 = {1{`RANDOM}};
  _T_6887_1153 = _RAND_1216[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1217 = {1{`RANDOM}};
  _T_6887_1154 = _RAND_1217[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1218 = {1{`RANDOM}};
  _T_6887_1155 = _RAND_1218[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1219 = {1{`RANDOM}};
  _T_6887_1156 = _RAND_1219[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1220 = {1{`RANDOM}};
  _T_6887_1157 = _RAND_1220[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1221 = {1{`RANDOM}};
  _T_6887_1158 = _RAND_1221[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1222 = {1{`RANDOM}};
  _T_6887_1159 = _RAND_1222[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1223 = {1{`RANDOM}};
  _T_6887_1160 = _RAND_1223[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1224 = {1{`RANDOM}};
  _T_6887_1161 = _RAND_1224[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1225 = {1{`RANDOM}};
  _T_6887_1162 = _RAND_1225[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1226 = {1{`RANDOM}};
  _T_6887_1163 = _RAND_1226[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1227 = {1{`RANDOM}};
  _T_6887_1164 = _RAND_1227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1228 = {1{`RANDOM}};
  _T_6887_1165 = _RAND_1228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1229 = {1{`RANDOM}};
  _T_6887_1166 = _RAND_1229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1230 = {1{`RANDOM}};
  _T_6887_1167 = _RAND_1230[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1231 = {1{`RANDOM}};
  _T_6887_1168 = _RAND_1231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1232 = {1{`RANDOM}};
  _T_6887_1169 = _RAND_1232[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1233 = {1{`RANDOM}};
  _T_6887_1170 = _RAND_1233[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1234 = {1{`RANDOM}};
  _T_6887_1171 = _RAND_1234[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1235 = {1{`RANDOM}};
  _T_6887_1172 = _RAND_1235[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1236 = {1{`RANDOM}};
  _T_6887_1173 = _RAND_1236[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1237 = {1{`RANDOM}};
  _T_6887_1174 = _RAND_1237[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1238 = {1{`RANDOM}};
  _T_6887_1175 = _RAND_1238[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1239 = {1{`RANDOM}};
  _T_6887_1176 = _RAND_1239[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1240 = {1{`RANDOM}};
  _T_6887_1177 = _RAND_1240[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1241 = {1{`RANDOM}};
  _T_6887_1178 = _RAND_1241[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1242 = {1{`RANDOM}};
  _T_6887_1179 = _RAND_1242[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1243 = {1{`RANDOM}};
  _T_6887_1180 = _RAND_1243[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1244 = {1{`RANDOM}};
  _T_6887_1181 = _RAND_1244[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1245 = {1{`RANDOM}};
  _T_6887_1182 = _RAND_1245[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1246 = {1{`RANDOM}};
  _T_6887_1183 = _RAND_1246[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1247 = {1{`RANDOM}};
  _T_6887_1184 = _RAND_1247[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1248 = {1{`RANDOM}};
  _T_6887_1185 = _RAND_1248[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1249 = {1{`RANDOM}};
  _T_6887_1186 = _RAND_1249[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1250 = {1{`RANDOM}};
  _T_6887_1187 = _RAND_1250[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1251 = {1{`RANDOM}};
  _T_6887_1188 = _RAND_1251[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1252 = {1{`RANDOM}};
  _T_6887_1189 = _RAND_1252[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1253 = {1{`RANDOM}};
  _T_6887_1190 = _RAND_1253[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1254 = {1{`RANDOM}};
  _T_6887_1191 = _RAND_1254[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1255 = {1{`RANDOM}};
  _T_6887_1192 = _RAND_1255[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1256 = {1{`RANDOM}};
  _T_6887_1193 = _RAND_1256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1257 = {1{`RANDOM}};
  _T_6887_1194 = _RAND_1257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1258 = {1{`RANDOM}};
  _T_6887_1195 = _RAND_1258[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1259 = {1{`RANDOM}};
  _T_6887_1196 = _RAND_1259[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1260 = {1{`RANDOM}};
  _T_6887_1197 = _RAND_1260[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1261 = {1{`RANDOM}};
  _T_6887_1198 = _RAND_1261[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1262 = {1{`RANDOM}};
  _T_6887_1199 = _RAND_1262[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1263 = {1{`RANDOM}};
  _T_6887_1200 = _RAND_1263[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1264 = {1{`RANDOM}};
  _T_6887_1201 = _RAND_1264[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1265 = {1{`RANDOM}};
  _T_6887_1202 = _RAND_1265[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1266 = {1{`RANDOM}};
  _T_6887_1203 = _RAND_1266[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1267 = {1{`RANDOM}};
  _T_6887_1204 = _RAND_1267[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1268 = {1{`RANDOM}};
  _T_6887_1205 = _RAND_1268[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1269 = {1{`RANDOM}};
  _T_6887_1206 = _RAND_1269[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1270 = {1{`RANDOM}};
  _T_6887_1207 = _RAND_1270[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1271 = {1{`RANDOM}};
  _T_6887_1208 = _RAND_1271[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1272 = {1{`RANDOM}};
  _T_6887_1209 = _RAND_1272[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1273 = {1{`RANDOM}};
  _T_6887_1210 = _RAND_1273[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1274 = {1{`RANDOM}};
  _T_6887_1211 = _RAND_1274[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1275 = {1{`RANDOM}};
  _T_6887_1212 = _RAND_1275[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1276 = {1{`RANDOM}};
  _T_6887_1213 = _RAND_1276[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1277 = {1{`RANDOM}};
  _T_6887_1214 = _RAND_1277[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1278 = {1{`RANDOM}};
  _T_6887_1215 = _RAND_1278[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1279 = {1{`RANDOM}};
  _T_6887_1216 = _RAND_1279[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1280 = {1{`RANDOM}};
  _T_6887_1217 = _RAND_1280[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1281 = {1{`RANDOM}};
  _T_6887_1218 = _RAND_1281[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1282 = {1{`RANDOM}};
  _T_6887_1219 = _RAND_1282[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1283 = {1{`RANDOM}};
  _T_6887_1220 = _RAND_1283[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1284 = {1{`RANDOM}};
  _T_6887_1221 = _RAND_1284[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1285 = {1{`RANDOM}};
  _T_6887_1222 = _RAND_1285[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1286 = {1{`RANDOM}};
  _T_6887_1223 = _RAND_1286[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1287 = {1{`RANDOM}};
  _T_6887_1224 = _RAND_1287[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1288 = {1{`RANDOM}};
  _T_6887_1225 = _RAND_1288[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1289 = {1{`RANDOM}};
  _T_6887_1226 = _RAND_1289[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1290 = {1{`RANDOM}};
  _T_6887_1227 = _RAND_1290[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1291 = {1{`RANDOM}};
  _T_6887_1228 = _RAND_1291[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1292 = {1{`RANDOM}};
  _T_6887_1229 = _RAND_1292[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1293 = {1{`RANDOM}};
  _T_6887_1230 = _RAND_1293[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1294 = {1{`RANDOM}};
  _T_6887_1231 = _RAND_1294[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1295 = {1{`RANDOM}};
  _T_6887_1232 = _RAND_1295[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1296 = {1{`RANDOM}};
  _T_6887_1233 = _RAND_1296[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1297 = {1{`RANDOM}};
  _T_6887_1234 = _RAND_1297[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1298 = {1{`RANDOM}};
  _T_6887_1235 = _RAND_1298[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1299 = {1{`RANDOM}};
  _T_6887_1236 = _RAND_1299[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1300 = {1{`RANDOM}};
  _T_6887_1237 = _RAND_1300[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1301 = {1{`RANDOM}};
  _T_6887_1238 = _RAND_1301[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1302 = {1{`RANDOM}};
  _T_6887_1239 = _RAND_1302[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1303 = {1{`RANDOM}};
  _T_6887_1240 = _RAND_1303[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1304 = {1{`RANDOM}};
  _T_6887_1241 = _RAND_1304[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1305 = {1{`RANDOM}};
  _T_6887_1242 = _RAND_1305[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1306 = {1{`RANDOM}};
  _T_6887_1243 = _RAND_1306[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1307 = {1{`RANDOM}};
  _T_6887_1244 = _RAND_1307[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1308 = {1{`RANDOM}};
  _T_6887_1245 = _RAND_1308[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1309 = {1{`RANDOM}};
  _T_6887_1246 = _RAND_1309[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1310 = {1{`RANDOM}};
  _T_6887_1247 = _RAND_1310[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1311 = {1{`RANDOM}};
  _T_6887_1248 = _RAND_1311[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1312 = {1{`RANDOM}};
  _T_6887_1249 = _RAND_1312[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1313 = {1{`RANDOM}};
  _T_6887_1250 = _RAND_1313[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1314 = {1{`RANDOM}};
  _T_6887_1251 = _RAND_1314[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1315 = {1{`RANDOM}};
  _T_6887_1252 = _RAND_1315[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1316 = {1{`RANDOM}};
  _T_6887_1253 = _RAND_1316[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1317 = {1{`RANDOM}};
  _T_6887_1254 = _RAND_1317[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1318 = {1{`RANDOM}};
  _T_6887_1255 = _RAND_1318[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1319 = {1{`RANDOM}};
  _T_6887_1256 = _RAND_1319[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1320 = {1{`RANDOM}};
  _T_6887_1257 = _RAND_1320[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1321 = {1{`RANDOM}};
  _T_6887_1258 = _RAND_1321[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1322 = {1{`RANDOM}};
  _T_6887_1259 = _RAND_1322[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1323 = {1{`RANDOM}};
  _T_6887_1260 = _RAND_1323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1324 = {1{`RANDOM}};
  _T_6887_1261 = _RAND_1324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1325 = {1{`RANDOM}};
  _T_6887_1262 = _RAND_1325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1326 = {1{`RANDOM}};
  _T_6887_1263 = _RAND_1326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1327 = {1{`RANDOM}};
  _T_6887_1264 = _RAND_1327[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1328 = {1{`RANDOM}};
  _T_6887_1265 = _RAND_1328[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1329 = {1{`RANDOM}};
  _T_6887_1266 = _RAND_1329[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1330 = {1{`RANDOM}};
  _T_6887_1267 = _RAND_1330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1331 = {1{`RANDOM}};
  _T_6887_1268 = _RAND_1331[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1332 = {1{`RANDOM}};
  _T_6887_1269 = _RAND_1332[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1333 = {1{`RANDOM}};
  _T_6887_1270 = _RAND_1333[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1334 = {1{`RANDOM}};
  _T_6887_1271 = _RAND_1334[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1335 = {1{`RANDOM}};
  _T_6887_1272 = _RAND_1335[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1336 = {1{`RANDOM}};
  _T_6887_1273 = _RAND_1336[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1337 = {1{`RANDOM}};
  _T_6887_1274 = _RAND_1337[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1338 = {1{`RANDOM}};
  _T_6887_1275 = _RAND_1338[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1339 = {1{`RANDOM}};
  _T_6887_1276 = _RAND_1339[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1340 = {1{`RANDOM}};
  _T_6887_1277 = _RAND_1340[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1341 = {1{`RANDOM}};
  _T_6887_1278 = _RAND_1341[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1342 = {1{`RANDOM}};
  _T_6887_1279 = _RAND_1342[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1343 = {1{`RANDOM}};
  _T_6887_1280 = _RAND_1343[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1344 = {1{`RANDOM}};
  _T_6887_1281 = _RAND_1344[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1345 = {1{`RANDOM}};
  _T_6887_1282 = _RAND_1345[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1346 = {1{`RANDOM}};
  _T_6887_1283 = _RAND_1346[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1347 = {1{`RANDOM}};
  _T_6887_1284 = _RAND_1347[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1348 = {1{`RANDOM}};
  _T_6887_1285 = _RAND_1348[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1349 = {1{`RANDOM}};
  _T_6887_1286 = _RAND_1349[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1350 = {1{`RANDOM}};
  _T_6887_1287 = _RAND_1350[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1351 = {1{`RANDOM}};
  _T_6887_1288 = _RAND_1351[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1352 = {1{`RANDOM}};
  _T_6887_1289 = _RAND_1352[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1353 = {1{`RANDOM}};
  _T_6887_1290 = _RAND_1353[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1354 = {1{`RANDOM}};
  _T_6887_1291 = _RAND_1354[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1355 = {1{`RANDOM}};
  _T_6887_1292 = _RAND_1355[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1356 = {1{`RANDOM}};
  _T_6887_1293 = _RAND_1356[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1357 = {1{`RANDOM}};
  _T_6887_1294 = _RAND_1357[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1358 = {1{`RANDOM}};
  _T_6887_1295 = _RAND_1358[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1359 = {1{`RANDOM}};
  _T_6887_1296 = _RAND_1359[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1360 = {1{`RANDOM}};
  _T_6887_1297 = _RAND_1360[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1361 = {1{`RANDOM}};
  _T_6887_1298 = _RAND_1361[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1362 = {1{`RANDOM}};
  _T_6887_1299 = _RAND_1362[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1363 = {1{`RANDOM}};
  _T_6887_1300 = _RAND_1363[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1364 = {1{`RANDOM}};
  _T_6887_1301 = _RAND_1364[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1365 = {1{`RANDOM}};
  _T_6887_1302 = _RAND_1365[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1366 = {1{`RANDOM}};
  _T_6887_1303 = _RAND_1366[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1367 = {1{`RANDOM}};
  _T_6887_1304 = _RAND_1367[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1368 = {1{`RANDOM}};
  _T_6887_1305 = _RAND_1368[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1369 = {1{`RANDOM}};
  _T_6887_1306 = _RAND_1369[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1370 = {1{`RANDOM}};
  _T_6887_1307 = _RAND_1370[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1371 = {1{`RANDOM}};
  _T_6887_1308 = _RAND_1371[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1372 = {1{`RANDOM}};
  _T_6887_1309 = _RAND_1372[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1373 = {1{`RANDOM}};
  _T_6887_1310 = _RAND_1373[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1374 = {1{`RANDOM}};
  _T_6887_1311 = _RAND_1374[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1375 = {1{`RANDOM}};
  _T_6887_1312 = _RAND_1375[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1376 = {1{`RANDOM}};
  _T_6887_1313 = _RAND_1376[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1377 = {1{`RANDOM}};
  _T_6887_1314 = _RAND_1377[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1378 = {1{`RANDOM}};
  _T_6887_1315 = _RAND_1378[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1379 = {1{`RANDOM}};
  _T_6887_1316 = _RAND_1379[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1380 = {1{`RANDOM}};
  _T_6887_1317 = _RAND_1380[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1381 = {1{`RANDOM}};
  _T_6887_1318 = _RAND_1381[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1382 = {1{`RANDOM}};
  _T_6887_1319 = _RAND_1382[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1383 = {1{`RANDOM}};
  _T_6887_1320 = _RAND_1383[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1384 = {1{`RANDOM}};
  _T_6887_1321 = _RAND_1384[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1385 = {1{`RANDOM}};
  _T_6887_1322 = _RAND_1385[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1386 = {1{`RANDOM}};
  _T_6887_1323 = _RAND_1386[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1387 = {1{`RANDOM}};
  _T_6887_1324 = _RAND_1387[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1388 = {1{`RANDOM}};
  _T_6887_1325 = _RAND_1388[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1389 = {1{`RANDOM}};
  _T_6887_1326 = _RAND_1389[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1390 = {1{`RANDOM}};
  _T_6887_1327 = _RAND_1390[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1391 = {1{`RANDOM}};
  _T_6887_1328 = _RAND_1391[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1392 = {1{`RANDOM}};
  _T_6887_1329 = _RAND_1392[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1393 = {1{`RANDOM}};
  _T_6887_1330 = _RAND_1393[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1394 = {1{`RANDOM}};
  _T_6887_1331 = _RAND_1394[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1395 = {1{`RANDOM}};
  _T_6887_1332 = _RAND_1395[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1396 = {1{`RANDOM}};
  _T_6887_1333 = _RAND_1396[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1397 = {1{`RANDOM}};
  _T_6887_1334 = _RAND_1397[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1398 = {1{`RANDOM}};
  _T_6887_1335 = _RAND_1398[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1399 = {1{`RANDOM}};
  _T_6887_1336 = _RAND_1399[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1400 = {1{`RANDOM}};
  _T_6887_1337 = _RAND_1400[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1401 = {1{`RANDOM}};
  _T_6887_1338 = _RAND_1401[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1402 = {1{`RANDOM}};
  _T_6887_1339 = _RAND_1402[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1403 = {1{`RANDOM}};
  _T_6887_1340 = _RAND_1403[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1404 = {1{`RANDOM}};
  _T_6887_1341 = _RAND_1404[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1405 = {1{`RANDOM}};
  _T_6887_1342 = _RAND_1405[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1406 = {1{`RANDOM}};
  _T_6887_1343 = _RAND_1406[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1407 = {1{`RANDOM}};
  _T_6887_1344 = _RAND_1407[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1408 = {1{`RANDOM}};
  _T_6887_1345 = _RAND_1408[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1409 = {1{`RANDOM}};
  _T_6887_1346 = _RAND_1409[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1410 = {1{`RANDOM}};
  _T_6887_1347 = _RAND_1410[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1411 = {1{`RANDOM}};
  _T_6887_1348 = _RAND_1411[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1412 = {1{`RANDOM}};
  _T_6887_1349 = _RAND_1412[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1413 = {1{`RANDOM}};
  _T_6887_1350 = _RAND_1413[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1414 = {1{`RANDOM}};
  _T_6887_1351 = _RAND_1414[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1415 = {1{`RANDOM}};
  _T_6887_1352 = _RAND_1415[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1416 = {1{`RANDOM}};
  _T_6887_1353 = _RAND_1416[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1417 = {1{`RANDOM}};
  _T_6887_1354 = _RAND_1417[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1418 = {1{`RANDOM}};
  _T_6887_1355 = _RAND_1418[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1419 = {1{`RANDOM}};
  _T_6887_1356 = _RAND_1419[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1420 = {1{`RANDOM}};
  _T_6887_1357 = _RAND_1420[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1421 = {1{`RANDOM}};
  _T_6887_1358 = _RAND_1421[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1422 = {1{`RANDOM}};
  _T_6887_1359 = _RAND_1422[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1423 = {1{`RANDOM}};
  _T_6887_1360 = _RAND_1423[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1424 = {1{`RANDOM}};
  _T_6887_1361 = _RAND_1424[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1425 = {1{`RANDOM}};
  _T_6887_1362 = _RAND_1425[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1426 = {1{`RANDOM}};
  _T_6887_1363 = _RAND_1426[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1427 = {1{`RANDOM}};
  _T_6887_1364 = _RAND_1427[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1428 = {1{`RANDOM}};
  _T_6887_1365 = _RAND_1428[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1429 = {1{`RANDOM}};
  _T_6887_1366 = _RAND_1429[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1430 = {1{`RANDOM}};
  _T_6887_1367 = _RAND_1430[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1431 = {1{`RANDOM}};
  _T_6887_1368 = _RAND_1431[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1432 = {1{`RANDOM}};
  _T_6887_1369 = _RAND_1432[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1433 = {1{`RANDOM}};
  _T_6887_1370 = _RAND_1433[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1434 = {1{`RANDOM}};
  _T_6887_1371 = _RAND_1434[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1435 = {1{`RANDOM}};
  _T_6887_1372 = _RAND_1435[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1436 = {1{`RANDOM}};
  _T_6887_1373 = _RAND_1436[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1437 = {1{`RANDOM}};
  _T_6887_1374 = _RAND_1437[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1438 = {1{`RANDOM}};
  _T_6887_1375 = _RAND_1438[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1439 = {1{`RANDOM}};
  _T_6887_1376 = _RAND_1439[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1440 = {1{`RANDOM}};
  _T_6887_1377 = _RAND_1440[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1441 = {1{`RANDOM}};
  _T_6887_1378 = _RAND_1441[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1442 = {1{`RANDOM}};
  _T_6887_1379 = _RAND_1442[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1443 = {1{`RANDOM}};
  _T_6887_1380 = _RAND_1443[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1444 = {1{`RANDOM}};
  _T_6887_1381 = _RAND_1444[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1445 = {1{`RANDOM}};
  _T_6887_1382 = _RAND_1445[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1446 = {1{`RANDOM}};
  _T_6887_1383 = _RAND_1446[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1447 = {1{`RANDOM}};
  _T_6887_1384 = _RAND_1447[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1448 = {1{`RANDOM}};
  _T_6887_1385 = _RAND_1448[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1449 = {1{`RANDOM}};
  _T_6887_1386 = _RAND_1449[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1450 = {1{`RANDOM}};
  _T_6887_1387 = _RAND_1450[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1451 = {1{`RANDOM}};
  _T_6887_1388 = _RAND_1451[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1452 = {1{`RANDOM}};
  _T_6887_1389 = _RAND_1452[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1453 = {1{`RANDOM}};
  _T_6887_1390 = _RAND_1453[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1454 = {1{`RANDOM}};
  _T_6887_1391 = _RAND_1454[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1455 = {1{`RANDOM}};
  _T_6887_1392 = _RAND_1455[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1456 = {1{`RANDOM}};
  _T_6887_1393 = _RAND_1456[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1457 = {1{`RANDOM}};
  _T_6887_1394 = _RAND_1457[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1458 = {1{`RANDOM}};
  _T_6887_1395 = _RAND_1458[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1459 = {1{`RANDOM}};
  _T_6887_1396 = _RAND_1459[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1460 = {1{`RANDOM}};
  _T_6887_1397 = _RAND_1460[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1461 = {1{`RANDOM}};
  _T_6887_1398 = _RAND_1461[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1462 = {1{`RANDOM}};
  _T_6887_1399 = _RAND_1462[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1463 = {1{`RANDOM}};
  _T_6887_1400 = _RAND_1463[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1464 = {1{`RANDOM}};
  _T_6887_1401 = _RAND_1464[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1465 = {1{`RANDOM}};
  _T_6887_1402 = _RAND_1465[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1466 = {1{`RANDOM}};
  _T_6887_1403 = _RAND_1466[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1467 = {1{`RANDOM}};
  _T_6887_1404 = _RAND_1467[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1468 = {1{`RANDOM}};
  _T_6887_1405 = _RAND_1468[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1469 = {1{`RANDOM}};
  _T_6887_1406 = _RAND_1469[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1470 = {1{`RANDOM}};
  _T_6887_1407 = _RAND_1470[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1471 = {1{`RANDOM}};
  _T_6887_1408 = _RAND_1471[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1472 = {1{`RANDOM}};
  _T_6887_1409 = _RAND_1472[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1473 = {1{`RANDOM}};
  _T_6887_1410 = _RAND_1473[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1474 = {1{`RANDOM}};
  _T_6887_1411 = _RAND_1474[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1475 = {1{`RANDOM}};
  _T_6887_1412 = _RAND_1475[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1476 = {1{`RANDOM}};
  _T_6887_1413 = _RAND_1476[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1477 = {1{`RANDOM}};
  _T_6887_1414 = _RAND_1477[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1478 = {1{`RANDOM}};
  _T_6887_1415 = _RAND_1478[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1479 = {1{`RANDOM}};
  _T_6887_1416 = _RAND_1479[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1480 = {1{`RANDOM}};
  _T_6887_1417 = _RAND_1480[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1481 = {1{`RANDOM}};
  _T_6887_1418 = _RAND_1481[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1482 = {1{`RANDOM}};
  _T_6887_1419 = _RAND_1482[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1483 = {1{`RANDOM}};
  _T_6887_1420 = _RAND_1483[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1484 = {1{`RANDOM}};
  _T_6887_1421 = _RAND_1484[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1485 = {1{`RANDOM}};
  _T_6887_1422 = _RAND_1485[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1486 = {1{`RANDOM}};
  _T_6887_1423 = _RAND_1486[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1487 = {1{`RANDOM}};
  _T_6887_1424 = _RAND_1487[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1488 = {1{`RANDOM}};
  _T_6887_1425 = _RAND_1488[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1489 = {1{`RANDOM}};
  _T_6887_1426 = _RAND_1489[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1490 = {1{`RANDOM}};
  _T_6887_1427 = _RAND_1490[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1491 = {1{`RANDOM}};
  _T_6887_1428 = _RAND_1491[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1492 = {1{`RANDOM}};
  _T_6887_1429 = _RAND_1492[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1493 = {1{`RANDOM}};
  _T_6887_1430 = _RAND_1493[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1494 = {1{`RANDOM}};
  _T_6887_1431 = _RAND_1494[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1495 = {1{`RANDOM}};
  _T_6887_1432 = _RAND_1495[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1496 = {1{`RANDOM}};
  _T_6887_1433 = _RAND_1496[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1497 = {1{`RANDOM}};
  _T_6887_1434 = _RAND_1497[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1498 = {1{`RANDOM}};
  _T_6887_1435 = _RAND_1498[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1499 = {1{`RANDOM}};
  _T_6887_1436 = _RAND_1499[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1500 = {1{`RANDOM}};
  _T_6887_1437 = _RAND_1500[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1501 = {1{`RANDOM}};
  _T_6887_1438 = _RAND_1501[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1502 = {1{`RANDOM}};
  _T_6887_1439 = _RAND_1502[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1503 = {1{`RANDOM}};
  _T_6887_1440 = _RAND_1503[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1504 = {1{`RANDOM}};
  _T_6887_1441 = _RAND_1504[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1505 = {1{`RANDOM}};
  _T_6887_1442 = _RAND_1505[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1506 = {1{`RANDOM}};
  _T_6887_1443 = _RAND_1506[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1507 = {1{`RANDOM}};
  _T_6887_1444 = _RAND_1507[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1508 = {1{`RANDOM}};
  _T_6887_1445 = _RAND_1508[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1509 = {1{`RANDOM}};
  _T_6887_1446 = _RAND_1509[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1510 = {1{`RANDOM}};
  _T_6887_1447 = _RAND_1510[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1511 = {1{`RANDOM}};
  _T_6887_1448 = _RAND_1511[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1512 = {1{`RANDOM}};
  _T_6887_1449 = _RAND_1512[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1513 = {1{`RANDOM}};
  _T_6887_1450 = _RAND_1513[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1514 = {1{`RANDOM}};
  _T_6887_1451 = _RAND_1514[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1515 = {1{`RANDOM}};
  _T_6887_1452 = _RAND_1515[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1516 = {1{`RANDOM}};
  _T_6887_1453 = _RAND_1516[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1517 = {1{`RANDOM}};
  _T_6887_1454 = _RAND_1517[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1518 = {1{`RANDOM}};
  _T_6887_1455 = _RAND_1518[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1519 = {1{`RANDOM}};
  _T_6887_1456 = _RAND_1519[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1520 = {1{`RANDOM}};
  _T_6887_1457 = _RAND_1520[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1521 = {1{`RANDOM}};
  _T_6887_1458 = _RAND_1521[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1522 = {1{`RANDOM}};
  _T_6887_1459 = _RAND_1522[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1523 = {1{`RANDOM}};
  _T_6887_1460 = _RAND_1523[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1524 = {1{`RANDOM}};
  _T_6887_1461 = _RAND_1524[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1525 = {1{`RANDOM}};
  _T_6887_1462 = _RAND_1525[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1526 = {1{`RANDOM}};
  _T_6887_1463 = _RAND_1526[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1527 = {1{`RANDOM}};
  _T_6887_1464 = _RAND_1527[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1528 = {1{`RANDOM}};
  _T_6887_1465 = _RAND_1528[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1529 = {1{`RANDOM}};
  _T_6887_1466 = _RAND_1529[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1530 = {1{`RANDOM}};
  _T_6887_1467 = _RAND_1530[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1531 = {1{`RANDOM}};
  _T_6887_1468 = _RAND_1531[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1532 = {1{`RANDOM}};
  _T_6887_1469 = _RAND_1532[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1533 = {1{`RANDOM}};
  _T_6887_1470 = _RAND_1533[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1534 = {1{`RANDOM}};
  _T_6887_1471 = _RAND_1534[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1535 = {1{`RANDOM}};
  _T_6887_1472 = _RAND_1535[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1536 = {1{`RANDOM}};
  _T_6887_1473 = _RAND_1536[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1537 = {1{`RANDOM}};
  _T_6887_1474 = _RAND_1537[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1538 = {1{`RANDOM}};
  _T_6887_1475 = _RAND_1538[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1539 = {1{`RANDOM}};
  _T_6887_1476 = _RAND_1539[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1540 = {1{`RANDOM}};
  _T_6887_1477 = _RAND_1540[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1541 = {1{`RANDOM}};
  _T_6887_1478 = _RAND_1541[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1542 = {1{`RANDOM}};
  _T_6887_1479 = _RAND_1542[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1543 = {1{`RANDOM}};
  _T_6887_1480 = _RAND_1543[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1544 = {1{`RANDOM}};
  _T_6887_1481 = _RAND_1544[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1545 = {1{`RANDOM}};
  _T_6887_1482 = _RAND_1545[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1546 = {1{`RANDOM}};
  _T_6887_1483 = _RAND_1546[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1547 = {1{`RANDOM}};
  _T_6887_1484 = _RAND_1547[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1548 = {1{`RANDOM}};
  _T_6887_1485 = _RAND_1548[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1549 = {1{`RANDOM}};
  _T_6887_1486 = _RAND_1549[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1550 = {1{`RANDOM}};
  _T_6887_1487 = _RAND_1550[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1551 = {1{`RANDOM}};
  _T_6887_1488 = _RAND_1551[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1552 = {1{`RANDOM}};
  _T_6887_1489 = _RAND_1552[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1553 = {1{`RANDOM}};
  _T_6887_1490 = _RAND_1553[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1554 = {1{`RANDOM}};
  _T_6887_1491 = _RAND_1554[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1555 = {1{`RANDOM}};
  _T_6887_1492 = _RAND_1555[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1556 = {1{`RANDOM}};
  _T_6887_1493 = _RAND_1556[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1557 = {1{`RANDOM}};
  _T_6887_1494 = _RAND_1557[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1558 = {1{`RANDOM}};
  _T_6887_1495 = _RAND_1558[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1559 = {1{`RANDOM}};
  _T_6887_1496 = _RAND_1559[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1560 = {1{`RANDOM}};
  _T_6887_1497 = _RAND_1560[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1561 = {1{`RANDOM}};
  _T_6887_1498 = _RAND_1561[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1562 = {1{`RANDOM}};
  _T_6887_1499 = _RAND_1562[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1563 = {1{`RANDOM}};
  _T_6887_1500 = _RAND_1563[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1564 = {1{`RANDOM}};
  _T_6887_1501 = _RAND_1564[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1565 = {1{`RANDOM}};
  _T_6887_1502 = _RAND_1565[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1566 = {1{`RANDOM}};
  _T_6887_1503 = _RAND_1566[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1567 = {1{`RANDOM}};
  _T_6887_1504 = _RAND_1567[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1568 = {1{`RANDOM}};
  _T_6887_1505 = _RAND_1568[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1569 = {1{`RANDOM}};
  _T_6887_1506 = _RAND_1569[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1570 = {1{`RANDOM}};
  _T_6887_1507 = _RAND_1570[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1571 = {1{`RANDOM}};
  _T_6887_1508 = _RAND_1571[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1572 = {1{`RANDOM}};
  _T_6887_1509 = _RAND_1572[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1573 = {1{`RANDOM}};
  _T_6887_1510 = _RAND_1573[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1574 = {1{`RANDOM}};
  _T_6887_1511 = _RAND_1574[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1575 = {1{`RANDOM}};
  _T_6887_1512 = _RAND_1575[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1576 = {1{`RANDOM}};
  _T_6887_1513 = _RAND_1576[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1577 = {1{`RANDOM}};
  _T_6887_1514 = _RAND_1577[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1578 = {1{`RANDOM}};
  _T_6887_1515 = _RAND_1578[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1579 = {1{`RANDOM}};
  _T_6887_1516 = _RAND_1579[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1580 = {1{`RANDOM}};
  _T_6887_1517 = _RAND_1580[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1581 = {1{`RANDOM}};
  _T_6887_1518 = _RAND_1581[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1582 = {1{`RANDOM}};
  _T_6887_1519 = _RAND_1582[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1583 = {1{`RANDOM}};
  _T_6887_1520 = _RAND_1583[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1584 = {1{`RANDOM}};
  _T_6887_1521 = _RAND_1584[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1585 = {1{`RANDOM}};
  _T_6887_1522 = _RAND_1585[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1586 = {1{`RANDOM}};
  _T_6887_1523 = _RAND_1586[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1587 = {1{`RANDOM}};
  _T_6887_1524 = _RAND_1587[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1588 = {1{`RANDOM}};
  _T_6887_1525 = _RAND_1588[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1589 = {1{`RANDOM}};
  _T_6887_1526 = _RAND_1589[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1590 = {1{`RANDOM}};
  _T_6887_1527 = _RAND_1590[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1591 = {1{`RANDOM}};
  _T_6887_1528 = _RAND_1591[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1592 = {1{`RANDOM}};
  _T_6887_1529 = _RAND_1592[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1593 = {1{`RANDOM}};
  _T_6887_1530 = _RAND_1593[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1594 = {1{`RANDOM}};
  _T_6887_1531 = _RAND_1594[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1595 = {1{`RANDOM}};
  _T_6887_1532 = _RAND_1595[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1596 = {1{`RANDOM}};
  _T_6887_1533 = _RAND_1596[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1597 = {1{`RANDOM}};
  _T_6887_1534 = _RAND_1597[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1598 = {1{`RANDOM}};
  _T_6887_1535 = _RAND_1598[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1599 = {1{`RANDOM}};
  _T_6887_1536 = _RAND_1599[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1600 = {1{`RANDOM}};
  _T_6887_1537 = _RAND_1600[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1601 = {1{`RANDOM}};
  _T_6887_1538 = _RAND_1601[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1602 = {1{`RANDOM}};
  _T_6887_1539 = _RAND_1602[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1603 = {1{`RANDOM}};
  _T_6887_1540 = _RAND_1603[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1604 = {1{`RANDOM}};
  _T_6887_1541 = _RAND_1604[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1605 = {1{`RANDOM}};
  _T_6887_1542 = _RAND_1605[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1606 = {1{`RANDOM}};
  _T_6887_1543 = _RAND_1606[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1607 = {1{`RANDOM}};
  _T_6887_1544 = _RAND_1607[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1608 = {1{`RANDOM}};
  _T_6887_1545 = _RAND_1608[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1609 = {1{`RANDOM}};
  _T_6887_1546 = _RAND_1609[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1610 = {1{`RANDOM}};
  _T_6887_1547 = _RAND_1610[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1611 = {1{`RANDOM}};
  _T_6887_1548 = _RAND_1611[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1612 = {1{`RANDOM}};
  _T_6887_1549 = _RAND_1612[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1613 = {1{`RANDOM}};
  _T_6887_1550 = _RAND_1613[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1614 = {1{`RANDOM}};
  _T_6887_1551 = _RAND_1614[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1615 = {1{`RANDOM}};
  _T_6887_1552 = _RAND_1615[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1616 = {1{`RANDOM}};
  _T_6887_1553 = _RAND_1616[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1617 = {1{`RANDOM}};
  _T_6887_1554 = _RAND_1617[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1618 = {1{`RANDOM}};
  _T_6887_1555 = _RAND_1618[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1619 = {1{`RANDOM}};
  _T_6887_1556 = _RAND_1619[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1620 = {1{`RANDOM}};
  _T_6887_1557 = _RAND_1620[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1621 = {1{`RANDOM}};
  _T_6887_1558 = _RAND_1621[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1622 = {1{`RANDOM}};
  _T_6887_1559 = _RAND_1622[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1623 = {1{`RANDOM}};
  _T_6887_1560 = _RAND_1623[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1624 = {1{`RANDOM}};
  _T_6887_1561 = _RAND_1624[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1625 = {1{`RANDOM}};
  _T_6887_1562 = _RAND_1625[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1626 = {1{`RANDOM}};
  _T_6887_1563 = _RAND_1626[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1627 = {1{`RANDOM}};
  _T_6887_1564 = _RAND_1627[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1628 = {1{`RANDOM}};
  _T_6887_1565 = _RAND_1628[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1629 = {1{`RANDOM}};
  _T_6887_1566 = _RAND_1629[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1630 = {1{`RANDOM}};
  _T_6887_1567 = _RAND_1630[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1631 = {1{`RANDOM}};
  _T_6887_1568 = _RAND_1631[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1632 = {1{`RANDOM}};
  _T_6887_1569 = _RAND_1632[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1633 = {1{`RANDOM}};
  _T_6887_1570 = _RAND_1633[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1634 = {1{`RANDOM}};
  _T_6887_1571 = _RAND_1634[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1635 = {1{`RANDOM}};
  _T_6887_1572 = _RAND_1635[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1636 = {1{`RANDOM}};
  _T_6887_1573 = _RAND_1636[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1637 = {1{`RANDOM}};
  _T_6887_1574 = _RAND_1637[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1638 = {1{`RANDOM}};
  _T_6887_1575 = _RAND_1638[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1639 = {1{`RANDOM}};
  _T_6887_1576 = _RAND_1639[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1640 = {1{`RANDOM}};
  _T_6887_1577 = _RAND_1640[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1641 = {1{`RANDOM}};
  _T_6887_1578 = _RAND_1641[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1642 = {1{`RANDOM}};
  _T_6887_1579 = _RAND_1642[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1643 = {1{`RANDOM}};
  _T_6887_1580 = _RAND_1643[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1644 = {1{`RANDOM}};
  _T_6887_1581 = _RAND_1644[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1645 = {1{`RANDOM}};
  _T_6887_1582 = _RAND_1645[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1646 = {1{`RANDOM}};
  _T_6887_1583 = _RAND_1646[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1647 = {1{`RANDOM}};
  _T_6887_1584 = _RAND_1647[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1648 = {1{`RANDOM}};
  _T_6887_1585 = _RAND_1648[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1649 = {1{`RANDOM}};
  _T_6887_1586 = _RAND_1649[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1650 = {1{`RANDOM}};
  _T_6887_1587 = _RAND_1650[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1651 = {1{`RANDOM}};
  _T_6887_1588 = _RAND_1651[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1652 = {1{`RANDOM}};
  _T_6887_1589 = _RAND_1652[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1653 = {1{`RANDOM}};
  _T_6887_1590 = _RAND_1653[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1654 = {1{`RANDOM}};
  _T_6887_1591 = _RAND_1654[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1655 = {1{`RANDOM}};
  _T_6887_1592 = _RAND_1655[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1656 = {1{`RANDOM}};
  _T_6887_1593 = _RAND_1656[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1657 = {1{`RANDOM}};
  _T_6887_1594 = _RAND_1657[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1658 = {1{`RANDOM}};
  _T_6887_1595 = _RAND_1658[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1659 = {1{`RANDOM}};
  _T_6887_1596 = _RAND_1659[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1660 = {1{`RANDOM}};
  _T_6887_1597 = _RAND_1660[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1661 = {1{`RANDOM}};
  _T_6887_1598 = _RAND_1661[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1662 = {1{`RANDOM}};
  _T_6887_1599 = _RAND_1662[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1663 = {1{`RANDOM}};
  _T_6887_1600 = _RAND_1663[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1664 = {1{`RANDOM}};
  _T_6887_1601 = _RAND_1664[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1665 = {1{`RANDOM}};
  _T_6887_1602 = _RAND_1665[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1666 = {1{`RANDOM}};
  _T_6887_1603 = _RAND_1666[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1667 = {1{`RANDOM}};
  _T_6887_1604 = _RAND_1667[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1668 = {1{`RANDOM}};
  _T_6887_1605 = _RAND_1668[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1669 = {1{`RANDOM}};
  _T_6887_1606 = _RAND_1669[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1670 = {1{`RANDOM}};
  _T_6887_1607 = _RAND_1670[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1671 = {1{`RANDOM}};
  _T_6887_1608 = _RAND_1671[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1672 = {1{`RANDOM}};
  _T_6887_1609 = _RAND_1672[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1673 = {1{`RANDOM}};
  _T_6887_1610 = _RAND_1673[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1674 = {1{`RANDOM}};
  _T_6887_1611 = _RAND_1674[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1675 = {1{`RANDOM}};
  _T_6887_1612 = _RAND_1675[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1676 = {1{`RANDOM}};
  _T_6887_1613 = _RAND_1676[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1677 = {1{`RANDOM}};
  _T_6887_1614 = _RAND_1677[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1678 = {1{`RANDOM}};
  _T_6887_1615 = _RAND_1678[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1679 = {1{`RANDOM}};
  _T_6887_1616 = _RAND_1679[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1680 = {1{`RANDOM}};
  _T_6887_1617 = _RAND_1680[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1681 = {1{`RANDOM}};
  _T_6887_1618 = _RAND_1681[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1682 = {1{`RANDOM}};
  _T_6887_1619 = _RAND_1682[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1683 = {1{`RANDOM}};
  _T_6887_1620 = _RAND_1683[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1684 = {1{`RANDOM}};
  _T_6887_1621 = _RAND_1684[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1685 = {1{`RANDOM}};
  _T_6887_1622 = _RAND_1685[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1686 = {1{`RANDOM}};
  _T_6887_1623 = _RAND_1686[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1687 = {1{`RANDOM}};
  _T_6887_1624 = _RAND_1687[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1688 = {1{`RANDOM}};
  _T_6887_1625 = _RAND_1688[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1689 = {1{`RANDOM}};
  _T_6887_1626 = _RAND_1689[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1690 = {1{`RANDOM}};
  _T_6887_1627 = _RAND_1690[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1691 = {1{`RANDOM}};
  _T_6887_1628 = _RAND_1691[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1692 = {1{`RANDOM}};
  _T_6887_1629 = _RAND_1692[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1693 = {1{`RANDOM}};
  _T_6887_1630 = _RAND_1693[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1694 = {1{`RANDOM}};
  _T_6887_1631 = _RAND_1694[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1695 = {1{`RANDOM}};
  _T_6887_1632 = _RAND_1695[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1696 = {1{`RANDOM}};
  _T_6887_1633 = _RAND_1696[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1697 = {1{`RANDOM}};
  _T_6887_1634 = _RAND_1697[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1698 = {1{`RANDOM}};
  _T_6887_1635 = _RAND_1698[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1699 = {1{`RANDOM}};
  _T_6887_1636 = _RAND_1699[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1700 = {1{`RANDOM}};
  _T_6887_1637 = _RAND_1700[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1701 = {1{`RANDOM}};
  _T_6887_1638 = _RAND_1701[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1702 = {1{`RANDOM}};
  _T_6887_1639 = _RAND_1702[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1703 = {1{`RANDOM}};
  _T_6887_1640 = _RAND_1703[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1704 = {1{`RANDOM}};
  _T_6887_1641 = _RAND_1704[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1705 = {1{`RANDOM}};
  _T_6887_1642 = _RAND_1705[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1706 = {1{`RANDOM}};
  _T_6887_1643 = _RAND_1706[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1707 = {1{`RANDOM}};
  _T_6887_1644 = _RAND_1707[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1708 = {1{`RANDOM}};
  _T_6887_1645 = _RAND_1708[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1709 = {1{`RANDOM}};
  _T_6887_1646 = _RAND_1709[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1710 = {1{`RANDOM}};
  _T_6887_1647 = _RAND_1710[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1711 = {1{`RANDOM}};
  _T_6887_1648 = _RAND_1711[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1712 = {1{`RANDOM}};
  _T_6887_1649 = _RAND_1712[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1713 = {1{`RANDOM}};
  _T_6887_1650 = _RAND_1713[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1714 = {1{`RANDOM}};
  _T_6887_1651 = _RAND_1714[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1715 = {1{`RANDOM}};
  _T_6887_1652 = _RAND_1715[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1716 = {1{`RANDOM}};
  _T_6887_1653 = _RAND_1716[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1717 = {1{`RANDOM}};
  _T_6887_1654 = _RAND_1717[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1718 = {1{`RANDOM}};
  _T_6887_1655 = _RAND_1718[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1719 = {1{`RANDOM}};
  _T_6887_1656 = _RAND_1719[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1720 = {1{`RANDOM}};
  _T_6887_1657 = _RAND_1720[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1721 = {1{`RANDOM}};
  _T_6887_1658 = _RAND_1721[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1722 = {1{`RANDOM}};
  _T_6887_1659 = _RAND_1722[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1723 = {1{`RANDOM}};
  _T_6887_1660 = _RAND_1723[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1724 = {1{`RANDOM}};
  _T_6887_1661 = _RAND_1724[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1725 = {1{`RANDOM}};
  _T_6887_1662 = _RAND_1725[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1726 = {1{`RANDOM}};
  _T_6887_1663 = _RAND_1726[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1727 = {1{`RANDOM}};
  _T_6887_1664 = _RAND_1727[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1728 = {1{`RANDOM}};
  _T_6887_1665 = _RAND_1728[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1729 = {1{`RANDOM}};
  _T_6887_1666 = _RAND_1729[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1730 = {1{`RANDOM}};
  _T_6887_1667 = _RAND_1730[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1731 = {1{`RANDOM}};
  _T_6887_1668 = _RAND_1731[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1732 = {1{`RANDOM}};
  _T_6887_1669 = _RAND_1732[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1733 = {1{`RANDOM}};
  _T_6887_1670 = _RAND_1733[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1734 = {1{`RANDOM}};
  _T_6887_1671 = _RAND_1734[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1735 = {1{`RANDOM}};
  _T_6887_1672 = _RAND_1735[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1736 = {1{`RANDOM}};
  _T_6887_1673 = _RAND_1736[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1737 = {1{`RANDOM}};
  _T_6887_1674 = _RAND_1737[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1738 = {1{`RANDOM}};
  _T_6887_1675 = _RAND_1738[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1739 = {1{`RANDOM}};
  _T_6887_1676 = _RAND_1739[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1740 = {1{`RANDOM}};
  _T_6887_1677 = _RAND_1740[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1741 = {1{`RANDOM}};
  _T_6887_1678 = _RAND_1741[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1742 = {1{`RANDOM}};
  _T_6887_1679 = _RAND_1742[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1743 = {1{`RANDOM}};
  _T_6887_1680 = _RAND_1743[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1744 = {1{`RANDOM}};
  _T_6887_1681 = _RAND_1744[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1745 = {1{`RANDOM}};
  _T_6887_1682 = _RAND_1745[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1746 = {1{`RANDOM}};
  _T_6887_1683 = _RAND_1746[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1747 = {1{`RANDOM}};
  _T_6887_1684 = _RAND_1747[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1748 = {1{`RANDOM}};
  _T_6887_1685 = _RAND_1748[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1749 = {1{`RANDOM}};
  _T_6887_1686 = _RAND_1749[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1750 = {1{`RANDOM}};
  _T_6887_1687 = _RAND_1750[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1751 = {1{`RANDOM}};
  _T_6887_1688 = _RAND_1751[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1752 = {1{`RANDOM}};
  _T_6887_1689 = _RAND_1752[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1753 = {1{`RANDOM}};
  _T_6887_1690 = _RAND_1753[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1754 = {1{`RANDOM}};
  _T_6887_1691 = _RAND_1754[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1755 = {1{`RANDOM}};
  _T_6887_1692 = _RAND_1755[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1756 = {1{`RANDOM}};
  _T_6887_1693 = _RAND_1756[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1757 = {1{`RANDOM}};
  _T_6887_1694 = _RAND_1757[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1758 = {1{`RANDOM}};
  _T_6887_1695 = _RAND_1758[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1759 = {1{`RANDOM}};
  _T_6887_1696 = _RAND_1759[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1760 = {1{`RANDOM}};
  _T_6887_1697 = _RAND_1760[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1761 = {1{`RANDOM}};
  _T_6887_1698 = _RAND_1761[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1762 = {1{`RANDOM}};
  _T_6887_1699 = _RAND_1762[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1763 = {1{`RANDOM}};
  _T_6887_1700 = _RAND_1763[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1764 = {1{`RANDOM}};
  _T_6887_1701 = _RAND_1764[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1765 = {1{`RANDOM}};
  _T_6887_1702 = _RAND_1765[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1766 = {1{`RANDOM}};
  _T_6887_1703 = _RAND_1766[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1767 = {1{`RANDOM}};
  _T_6887_1704 = _RAND_1767[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1768 = {1{`RANDOM}};
  _T_6887_1705 = _RAND_1768[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1769 = {1{`RANDOM}};
  _T_6887_1706 = _RAND_1769[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1770 = {1{`RANDOM}};
  _T_6887_1707 = _RAND_1770[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1771 = {1{`RANDOM}};
  _T_6887_1708 = _RAND_1771[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1772 = {1{`RANDOM}};
  _T_6887_1709 = _RAND_1772[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1773 = {1{`RANDOM}};
  _T_6887_1710 = _RAND_1773[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1774 = {1{`RANDOM}};
  _T_6887_1711 = _RAND_1774[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1775 = {1{`RANDOM}};
  _T_6887_1712 = _RAND_1775[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1776 = {1{`RANDOM}};
  _T_6887_1713 = _RAND_1776[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1777 = {1{`RANDOM}};
  _T_6887_1714 = _RAND_1777[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1778 = {1{`RANDOM}};
  _T_6887_1715 = _RAND_1778[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1779 = {1{`RANDOM}};
  _T_6887_1716 = _RAND_1779[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1780 = {1{`RANDOM}};
  _T_6887_1717 = _RAND_1780[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1781 = {1{`RANDOM}};
  _T_6887_1718 = _RAND_1781[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1782 = {1{`RANDOM}};
  _T_6887_1719 = _RAND_1782[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1783 = {1{`RANDOM}};
  _T_6887_1720 = _RAND_1783[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1784 = {1{`RANDOM}};
  _T_6887_1721 = _RAND_1784[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1785 = {1{`RANDOM}};
  _T_6887_1722 = _RAND_1785[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1786 = {1{`RANDOM}};
  _T_6887_1723 = _RAND_1786[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1787 = {1{`RANDOM}};
  _T_6887_1724 = _RAND_1787[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1788 = {1{`RANDOM}};
  _T_6887_1725 = _RAND_1788[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1789 = {1{`RANDOM}};
  _T_6887_1726 = _RAND_1789[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1790 = {1{`RANDOM}};
  _T_6887_1727 = _RAND_1790[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1791 = {1{`RANDOM}};
  _T_6887_1728 = _RAND_1791[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1792 = {1{`RANDOM}};
  _T_6887_1729 = _RAND_1792[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1793 = {1{`RANDOM}};
  _T_6887_1730 = _RAND_1793[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1794 = {1{`RANDOM}};
  _T_6887_1731 = _RAND_1794[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1795 = {1{`RANDOM}};
  _T_6887_1732 = _RAND_1795[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1796 = {1{`RANDOM}};
  _T_6887_1733 = _RAND_1796[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1797 = {1{`RANDOM}};
  _T_6887_1734 = _RAND_1797[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1798 = {1{`RANDOM}};
  _T_6887_1735 = _RAND_1798[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1799 = {1{`RANDOM}};
  _T_6887_1736 = _RAND_1799[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1800 = {1{`RANDOM}};
  _T_6887_1737 = _RAND_1800[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1801 = {1{`RANDOM}};
  _T_6887_1738 = _RAND_1801[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1802 = {1{`RANDOM}};
  _T_6887_1739 = _RAND_1802[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1803 = {1{`RANDOM}};
  _T_6887_1740 = _RAND_1803[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1804 = {1{`RANDOM}};
  _T_6887_1741 = _RAND_1804[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1805 = {1{`RANDOM}};
  _T_6887_1742 = _RAND_1805[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1806 = {1{`RANDOM}};
  _T_6887_1743 = _RAND_1806[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1807 = {1{`RANDOM}};
  _T_6887_1744 = _RAND_1807[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1808 = {1{`RANDOM}};
  _T_6887_1745 = _RAND_1808[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1809 = {1{`RANDOM}};
  _T_6887_1746 = _RAND_1809[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1810 = {1{`RANDOM}};
  _T_6887_1747 = _RAND_1810[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1811 = {1{`RANDOM}};
  _T_6887_1748 = _RAND_1811[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1812 = {1{`RANDOM}};
  _T_6887_1749 = _RAND_1812[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1813 = {1{`RANDOM}};
  _T_6887_1750 = _RAND_1813[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1814 = {1{`RANDOM}};
  _T_6887_1751 = _RAND_1814[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1815 = {1{`RANDOM}};
  _T_6887_1752 = _RAND_1815[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1816 = {1{`RANDOM}};
  _T_6887_1753 = _RAND_1816[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1817 = {1{`RANDOM}};
  _T_6887_1754 = _RAND_1817[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1818 = {1{`RANDOM}};
  _T_6887_1755 = _RAND_1818[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1819 = {1{`RANDOM}};
  _T_6887_1756 = _RAND_1819[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1820 = {1{`RANDOM}};
  _T_6887_1757 = _RAND_1820[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1821 = {1{`RANDOM}};
  _T_6887_1758 = _RAND_1821[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1822 = {1{`RANDOM}};
  _T_6887_1759 = _RAND_1822[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1823 = {1{`RANDOM}};
  _T_6887_1760 = _RAND_1823[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1824 = {1{`RANDOM}};
  _T_6887_1761 = _RAND_1824[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1825 = {1{`RANDOM}};
  _T_6887_1762 = _RAND_1825[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1826 = {1{`RANDOM}};
  _T_6887_1763 = _RAND_1826[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1827 = {1{`RANDOM}};
  _T_6887_1764 = _RAND_1827[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1828 = {1{`RANDOM}};
  _T_6887_1765 = _RAND_1828[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1829 = {1{`RANDOM}};
  _T_6887_1766 = _RAND_1829[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1830 = {1{`RANDOM}};
  _T_6887_1767 = _RAND_1830[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1831 = {1{`RANDOM}};
  _T_6887_1768 = _RAND_1831[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1832 = {1{`RANDOM}};
  _T_6887_1769 = _RAND_1832[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1833 = {1{`RANDOM}};
  _T_6887_1770 = _RAND_1833[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1834 = {1{`RANDOM}};
  _T_6887_1771 = _RAND_1834[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1835 = {1{`RANDOM}};
  _T_6887_1772 = _RAND_1835[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1836 = {1{`RANDOM}};
  _T_6887_1773 = _RAND_1836[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1837 = {1{`RANDOM}};
  _T_6887_1774 = _RAND_1837[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1838 = {1{`RANDOM}};
  _T_6887_1775 = _RAND_1838[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1839 = {1{`RANDOM}};
  _T_6887_1776 = _RAND_1839[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1840 = {1{`RANDOM}};
  _T_6887_1777 = _RAND_1840[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1841 = {1{`RANDOM}};
  _T_6887_1778 = _RAND_1841[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1842 = {1{`RANDOM}};
  _T_6887_1779 = _RAND_1842[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1843 = {1{`RANDOM}};
  _T_6887_1780 = _RAND_1843[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1844 = {1{`RANDOM}};
  _T_6887_1781 = _RAND_1844[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1845 = {1{`RANDOM}};
  _T_6887_1782 = _RAND_1845[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1846 = {1{`RANDOM}};
  _T_6887_1783 = _RAND_1846[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1847 = {1{`RANDOM}};
  _T_6887_1784 = _RAND_1847[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1848 = {1{`RANDOM}};
  _T_6887_1785 = _RAND_1848[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1849 = {1{`RANDOM}};
  _T_6887_1786 = _RAND_1849[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1850 = {1{`RANDOM}};
  _T_6887_1787 = _RAND_1850[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1851 = {1{`RANDOM}};
  _T_6887_1788 = _RAND_1851[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1852 = {1{`RANDOM}};
  _T_6887_1789 = _RAND_1852[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1853 = {1{`RANDOM}};
  _T_6887_1790 = _RAND_1853[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1854 = {1{`RANDOM}};
  _T_6887_1791 = _RAND_1854[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1855 = {1{`RANDOM}};
  _T_6887_1792 = _RAND_1855[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1856 = {1{`RANDOM}};
  _T_6887_1793 = _RAND_1856[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1857 = {1{`RANDOM}};
  _T_6887_1794 = _RAND_1857[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1858 = {1{`RANDOM}};
  _T_6887_1795 = _RAND_1858[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1859 = {1{`RANDOM}};
  _T_6887_1796 = _RAND_1859[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1860 = {1{`RANDOM}};
  _T_6887_1797 = _RAND_1860[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1861 = {1{`RANDOM}};
  _T_6887_1798 = _RAND_1861[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1862 = {1{`RANDOM}};
  _T_6887_1799 = _RAND_1862[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1863 = {1{`RANDOM}};
  _T_6887_1800 = _RAND_1863[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1864 = {1{`RANDOM}};
  _T_6887_1801 = _RAND_1864[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1865 = {1{`RANDOM}};
  _T_6887_1802 = _RAND_1865[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1866 = {1{`RANDOM}};
  _T_6887_1803 = _RAND_1866[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1867 = {1{`RANDOM}};
  _T_6887_1804 = _RAND_1867[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1868 = {1{`RANDOM}};
  _T_6887_1805 = _RAND_1868[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1869 = {1{`RANDOM}};
  _T_6887_1806 = _RAND_1869[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1870 = {1{`RANDOM}};
  _T_6887_1807 = _RAND_1870[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1871 = {1{`RANDOM}};
  _T_6887_1808 = _RAND_1871[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1872 = {1{`RANDOM}};
  _T_6887_1809 = _RAND_1872[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1873 = {1{`RANDOM}};
  _T_6887_1810 = _RAND_1873[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1874 = {1{`RANDOM}};
  _T_6887_1811 = _RAND_1874[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1875 = {1{`RANDOM}};
  _T_6887_1812 = _RAND_1875[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1876 = {1{`RANDOM}};
  _T_6887_1813 = _RAND_1876[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1877 = {1{`RANDOM}};
  _T_6887_1814 = _RAND_1877[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1878 = {1{`RANDOM}};
  _T_6887_1815 = _RAND_1878[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1879 = {1{`RANDOM}};
  _T_6887_1816 = _RAND_1879[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1880 = {1{`RANDOM}};
  _T_6887_1817 = _RAND_1880[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1881 = {1{`RANDOM}};
  _T_6887_1818 = _RAND_1881[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1882 = {1{`RANDOM}};
  _T_6887_1819 = _RAND_1882[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1883 = {1{`RANDOM}};
  _T_6887_1820 = _RAND_1883[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1884 = {1{`RANDOM}};
  _T_6887_1821 = _RAND_1884[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1885 = {1{`RANDOM}};
  _T_6887_1822 = _RAND_1885[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1886 = {1{`RANDOM}};
  _T_6887_1823 = _RAND_1886[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1887 = {1{`RANDOM}};
  _T_6887_1824 = _RAND_1887[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1888 = {1{`RANDOM}};
  _T_6887_1825 = _RAND_1888[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1889 = {1{`RANDOM}};
  _T_6887_1826 = _RAND_1889[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1890 = {1{`RANDOM}};
  _T_6887_1827 = _RAND_1890[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1891 = {1{`RANDOM}};
  _T_6887_1828 = _RAND_1891[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1892 = {1{`RANDOM}};
  _T_6887_1829 = _RAND_1892[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1893 = {1{`RANDOM}};
  _T_6887_1830 = _RAND_1893[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1894 = {1{`RANDOM}};
  _T_6887_1831 = _RAND_1894[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1895 = {1{`RANDOM}};
  _T_6887_1832 = _RAND_1895[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1896 = {1{`RANDOM}};
  _T_6887_1833 = _RAND_1896[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1897 = {1{`RANDOM}};
  _T_6887_1834 = _RAND_1897[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1898 = {1{`RANDOM}};
  _T_6887_1835 = _RAND_1898[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1899 = {1{`RANDOM}};
  _T_6887_1836 = _RAND_1899[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1900 = {1{`RANDOM}};
  _T_6887_1837 = _RAND_1900[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1901 = {1{`RANDOM}};
  _T_6887_1838 = _RAND_1901[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1902 = {1{`RANDOM}};
  _T_6887_1839 = _RAND_1902[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1903 = {1{`RANDOM}};
  _T_6887_1840 = _RAND_1903[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1904 = {1{`RANDOM}};
  _T_6887_1841 = _RAND_1904[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1905 = {1{`RANDOM}};
  _T_6887_1842 = _RAND_1905[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1906 = {1{`RANDOM}};
  _T_6887_1843 = _RAND_1906[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1907 = {1{`RANDOM}};
  _T_6887_1844 = _RAND_1907[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1908 = {1{`RANDOM}};
  _T_6887_1845 = _RAND_1908[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1909 = {1{`RANDOM}};
  _T_6887_1846 = _RAND_1909[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1910 = {1{`RANDOM}};
  _T_6887_1847 = _RAND_1910[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1911 = {1{`RANDOM}};
  _T_6887_1848 = _RAND_1911[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1912 = {1{`RANDOM}};
  _T_6887_1849 = _RAND_1912[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1913 = {1{`RANDOM}};
  _T_6887_1850 = _RAND_1913[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1914 = {1{`RANDOM}};
  _T_6887_1851 = _RAND_1914[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1915 = {1{`RANDOM}};
  _T_6887_1852 = _RAND_1915[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1916 = {1{`RANDOM}};
  _T_6887_1853 = _RAND_1916[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1917 = {1{`RANDOM}};
  _T_6887_1854 = _RAND_1917[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1918 = {1{`RANDOM}};
  _T_6887_1855 = _RAND_1918[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1919 = {1{`RANDOM}};
  _T_6887_1856 = _RAND_1919[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1920 = {1{`RANDOM}};
  _T_6887_1857 = _RAND_1920[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1921 = {1{`RANDOM}};
  _T_6887_1858 = _RAND_1921[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1922 = {1{`RANDOM}};
  _T_6887_1859 = _RAND_1922[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1923 = {1{`RANDOM}};
  _T_6887_1860 = _RAND_1923[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1924 = {1{`RANDOM}};
  _T_6887_1861 = _RAND_1924[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1925 = {1{`RANDOM}};
  _T_6887_1862 = _RAND_1925[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1926 = {1{`RANDOM}};
  _T_6887_1863 = _RAND_1926[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1927 = {1{`RANDOM}};
  _T_6887_1864 = _RAND_1927[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1928 = {1{`RANDOM}};
  _T_6887_1865 = _RAND_1928[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1929 = {1{`RANDOM}};
  _T_6887_1866 = _RAND_1929[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1930 = {1{`RANDOM}};
  _T_6887_1867 = _RAND_1930[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1931 = {1{`RANDOM}};
  _T_6887_1868 = _RAND_1931[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1932 = {1{`RANDOM}};
  _T_6887_1869 = _RAND_1932[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1933 = {1{`RANDOM}};
  _T_6887_1870 = _RAND_1933[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1934 = {1{`RANDOM}};
  _T_6887_1871 = _RAND_1934[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1935 = {1{`RANDOM}};
  _T_6887_1872 = _RAND_1935[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1936 = {1{`RANDOM}};
  _T_6887_1873 = _RAND_1936[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1937 = {1{`RANDOM}};
  _T_6887_1874 = _RAND_1937[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1938 = {1{`RANDOM}};
  _T_6887_1875 = _RAND_1938[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1939 = {1{`RANDOM}};
  _T_6887_1876 = _RAND_1939[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1940 = {1{`RANDOM}};
  _T_6887_1877 = _RAND_1940[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1941 = {1{`RANDOM}};
  _T_6887_1878 = _RAND_1941[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1942 = {1{`RANDOM}};
  _T_6887_1879 = _RAND_1942[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1943 = {1{`RANDOM}};
  _T_6887_1880 = _RAND_1943[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1944 = {1{`RANDOM}};
  _T_6887_1881 = _RAND_1944[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1945 = {1{`RANDOM}};
  _T_6887_1882 = _RAND_1945[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1946 = {1{`RANDOM}};
  _T_6887_1883 = _RAND_1946[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1947 = {1{`RANDOM}};
  _T_6887_1884 = _RAND_1947[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1948 = {1{`RANDOM}};
  _T_6887_1885 = _RAND_1948[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1949 = {1{`RANDOM}};
  _T_6887_1886 = _RAND_1949[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1950 = {1{`RANDOM}};
  _T_6887_1887 = _RAND_1950[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1951 = {1{`RANDOM}};
  _T_6887_1888 = _RAND_1951[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1952 = {1{`RANDOM}};
  _T_6887_1889 = _RAND_1952[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1953 = {1{`RANDOM}};
  _T_6887_1890 = _RAND_1953[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1954 = {1{`RANDOM}};
  _T_6887_1891 = _RAND_1954[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1955 = {1{`RANDOM}};
  _T_6887_1892 = _RAND_1955[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1956 = {1{`RANDOM}};
  _T_6887_1893 = _RAND_1956[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1957 = {1{`RANDOM}};
  _T_6887_1894 = _RAND_1957[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1958 = {1{`RANDOM}};
  _T_6887_1895 = _RAND_1958[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1959 = {1{`RANDOM}};
  _T_6887_1896 = _RAND_1959[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1960 = {1{`RANDOM}};
  _T_6887_1897 = _RAND_1960[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1961 = {1{`RANDOM}};
  _T_6887_1898 = _RAND_1961[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1962 = {1{`RANDOM}};
  _T_6887_1899 = _RAND_1962[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1963 = {1{`RANDOM}};
  _T_6887_1900 = _RAND_1963[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1964 = {1{`RANDOM}};
  _T_6887_1901 = _RAND_1964[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1965 = {1{`RANDOM}};
  _T_6887_1902 = _RAND_1965[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1966 = {1{`RANDOM}};
  _T_6887_1903 = _RAND_1966[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1967 = {1{`RANDOM}};
  _T_6887_1904 = _RAND_1967[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1968 = {1{`RANDOM}};
  _T_6887_1905 = _RAND_1968[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1969 = {1{`RANDOM}};
  _T_6887_1906 = _RAND_1969[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1970 = {1{`RANDOM}};
  _T_6887_1907 = _RAND_1970[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1971 = {1{`RANDOM}};
  _T_6887_1908 = _RAND_1971[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1972 = {1{`RANDOM}};
  _T_6887_1909 = _RAND_1972[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1973 = {1{`RANDOM}};
  _T_6887_1910 = _RAND_1973[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1974 = {1{`RANDOM}};
  _T_6887_1911 = _RAND_1974[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1975 = {1{`RANDOM}};
  _T_6887_1912 = _RAND_1975[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1976 = {1{`RANDOM}};
  _T_6887_1913 = _RAND_1976[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1977 = {1{`RANDOM}};
  _T_6887_1914 = _RAND_1977[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1978 = {1{`RANDOM}};
  _T_6887_1915 = _RAND_1978[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1979 = {1{`RANDOM}};
  _T_6887_1916 = _RAND_1979[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1980 = {1{`RANDOM}};
  _T_6887_1917 = _RAND_1980[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1981 = {1{`RANDOM}};
  _T_6887_1918 = _RAND_1981[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1982 = {1{`RANDOM}};
  _T_6887_1919 = _RAND_1982[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1983 = {1{`RANDOM}};
  _T_6887_1920 = _RAND_1983[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1984 = {1{`RANDOM}};
  _T_6887_1921 = _RAND_1984[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1985 = {1{`RANDOM}};
  _T_6887_1922 = _RAND_1985[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1986 = {1{`RANDOM}};
  _T_6887_1923 = _RAND_1986[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1987 = {1{`RANDOM}};
  _T_6887_1924 = _RAND_1987[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1988 = {1{`RANDOM}};
  _T_6887_1925 = _RAND_1988[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1989 = {1{`RANDOM}};
  _T_6887_1926 = _RAND_1989[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1990 = {1{`RANDOM}};
  _T_6887_1927 = _RAND_1990[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1991 = {1{`RANDOM}};
  _T_6887_1928 = _RAND_1991[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1992 = {1{`RANDOM}};
  _T_6887_1929 = _RAND_1992[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1993 = {1{`RANDOM}};
  _T_6887_1930 = _RAND_1993[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1994 = {1{`RANDOM}};
  _T_6887_1931 = _RAND_1994[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1995 = {1{`RANDOM}};
  _T_6887_1932 = _RAND_1995[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1996 = {1{`RANDOM}};
  _T_6887_1933 = _RAND_1996[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1997 = {1{`RANDOM}};
  _T_6887_1934 = _RAND_1997[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1998 = {1{`RANDOM}};
  _T_6887_1935 = _RAND_1998[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1999 = {1{`RANDOM}};
  _T_6887_1936 = _RAND_1999[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2000 = {1{`RANDOM}};
  _T_6887_1937 = _RAND_2000[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2001 = {1{`RANDOM}};
  _T_6887_1938 = _RAND_2001[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2002 = {1{`RANDOM}};
  _T_6887_1939 = _RAND_2002[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2003 = {1{`RANDOM}};
  _T_6887_1940 = _RAND_2003[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2004 = {1{`RANDOM}};
  _T_6887_1941 = _RAND_2004[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2005 = {1{`RANDOM}};
  _T_6887_1942 = _RAND_2005[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2006 = {1{`RANDOM}};
  _T_6887_1943 = _RAND_2006[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2007 = {1{`RANDOM}};
  _T_6887_1944 = _RAND_2007[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2008 = {1{`RANDOM}};
  _T_6887_1945 = _RAND_2008[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2009 = {1{`RANDOM}};
  _T_6887_1946 = _RAND_2009[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2010 = {1{`RANDOM}};
  _T_6887_1947 = _RAND_2010[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2011 = {1{`RANDOM}};
  _T_6887_1948 = _RAND_2011[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2012 = {1{`RANDOM}};
  _T_6887_1949 = _RAND_2012[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2013 = {1{`RANDOM}};
  _T_6887_1950 = _RAND_2013[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2014 = {1{`RANDOM}};
  _T_6887_1951 = _RAND_2014[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2015 = {1{`RANDOM}};
  _T_6887_1952 = _RAND_2015[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2016 = {1{`RANDOM}};
  _T_6887_1953 = _RAND_2016[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2017 = {1{`RANDOM}};
  _T_6887_1954 = _RAND_2017[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2018 = {1{`RANDOM}};
  _T_6887_1955 = _RAND_2018[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2019 = {1{`RANDOM}};
  _T_6887_1956 = _RAND_2019[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2020 = {1{`RANDOM}};
  _T_6887_1957 = _RAND_2020[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2021 = {1{`RANDOM}};
  _T_6887_1958 = _RAND_2021[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2022 = {1{`RANDOM}};
  _T_6887_1959 = _RAND_2022[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2023 = {1{`RANDOM}};
  _T_6887_1960 = _RAND_2023[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2024 = {1{`RANDOM}};
  _T_6887_1961 = _RAND_2024[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2025 = {1{`RANDOM}};
  _T_6887_1962 = _RAND_2025[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2026 = {1{`RANDOM}};
  _T_6887_1963 = _RAND_2026[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2027 = {1{`RANDOM}};
  _T_6887_1964 = _RAND_2027[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2028 = {1{`RANDOM}};
  _T_6887_1965 = _RAND_2028[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2029 = {1{`RANDOM}};
  _T_6887_1966 = _RAND_2029[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2030 = {1{`RANDOM}};
  _T_6887_1967 = _RAND_2030[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2031 = {1{`RANDOM}};
  _T_6887_1968 = _RAND_2031[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2032 = {1{`RANDOM}};
  _T_6887_1969 = _RAND_2032[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2033 = {1{`RANDOM}};
  _T_6887_1970 = _RAND_2033[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2034 = {1{`RANDOM}};
  _T_6887_1971 = _RAND_2034[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2035 = {1{`RANDOM}};
  _T_6887_1972 = _RAND_2035[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2036 = {1{`RANDOM}};
  _T_6887_1973 = _RAND_2036[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2037 = {1{`RANDOM}};
  _T_6887_1974 = _RAND_2037[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2038 = {1{`RANDOM}};
  _T_6887_1975 = _RAND_2038[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2039 = {1{`RANDOM}};
  _T_6887_1976 = _RAND_2039[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2040 = {1{`RANDOM}};
  _T_6887_1977 = _RAND_2040[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2041 = {1{`RANDOM}};
  _T_6887_1978 = _RAND_2041[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2042 = {1{`RANDOM}};
  _T_6887_1979 = _RAND_2042[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2043 = {1{`RANDOM}};
  _T_6887_1980 = _RAND_2043[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2044 = {1{`RANDOM}};
  _T_6887_1981 = _RAND_2044[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2045 = {1{`RANDOM}};
  _T_6887_1982 = _RAND_2045[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2046 = {1{`RANDOM}};
  _T_6887_1983 = _RAND_2046[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2047 = {1{`RANDOM}};
  _T_6887_1984 = _RAND_2047[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2048 = {1{`RANDOM}};
  _T_6887_1985 = _RAND_2048[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2049 = {1{`RANDOM}};
  _T_6887_1986 = _RAND_2049[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2050 = {1{`RANDOM}};
  _T_6887_1987 = _RAND_2050[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2051 = {1{`RANDOM}};
  _T_6887_1988 = _RAND_2051[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2052 = {1{`RANDOM}};
  _T_6887_1989 = _RAND_2052[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2053 = {1{`RANDOM}};
  _T_6887_1990 = _RAND_2053[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2054 = {1{`RANDOM}};
  _T_6887_1991 = _RAND_2054[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2055 = {1{`RANDOM}};
  _T_6887_1992 = _RAND_2055[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2056 = {1{`RANDOM}};
  _T_6887_1993 = _RAND_2056[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2057 = {1{`RANDOM}};
  _T_6887_1994 = _RAND_2057[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2058 = {1{`RANDOM}};
  _T_6887_1995 = _RAND_2058[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2059 = {1{`RANDOM}};
  _T_6887_1996 = _RAND_2059[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2060 = {1{`RANDOM}};
  _T_6887_1997 = _RAND_2060[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2061 = {1{`RANDOM}};
  _T_6887_1998 = _RAND_2061[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2062 = {1{`RANDOM}};
  _T_6887_1999 = _RAND_2062[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2063 = {1{`RANDOM}};
  _T_6887_2000 = _RAND_2063[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2064 = {1{`RANDOM}};
  _T_6887_2001 = _RAND_2064[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2065 = {1{`RANDOM}};
  _T_6887_2002 = _RAND_2065[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2066 = {1{`RANDOM}};
  _T_6887_2003 = _RAND_2066[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2067 = {1{`RANDOM}};
  _T_6887_2004 = _RAND_2067[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2068 = {1{`RANDOM}};
  _T_6887_2005 = _RAND_2068[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2069 = {1{`RANDOM}};
  _T_6887_2006 = _RAND_2069[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2070 = {1{`RANDOM}};
  _T_6887_2007 = _RAND_2070[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2071 = {1{`RANDOM}};
  _T_6887_2008 = _RAND_2071[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2072 = {1{`RANDOM}};
  _T_6887_2009 = _RAND_2072[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2073 = {1{`RANDOM}};
  _T_6887_2010 = _RAND_2073[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2074 = {1{`RANDOM}};
  _T_6887_2011 = _RAND_2074[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2075 = {1{`RANDOM}};
  _T_6887_2012 = _RAND_2075[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2076 = {1{`RANDOM}};
  _T_6887_2013 = _RAND_2076[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2077 = {1{`RANDOM}};
  _T_6887_2014 = _RAND_2077[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2078 = {1{`RANDOM}};
  _T_6887_2015 = _RAND_2078[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2079 = {1{`RANDOM}};
  _T_6887_2016 = _RAND_2079[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2080 = {1{`RANDOM}};
  _T_6887_2017 = _RAND_2080[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2081 = {1{`RANDOM}};
  _T_6887_2018 = _RAND_2081[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2082 = {1{`RANDOM}};
  _T_6887_2019 = _RAND_2082[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2083 = {1{`RANDOM}};
  _T_6887_2020 = _RAND_2083[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2084 = {1{`RANDOM}};
  _T_6887_2021 = _RAND_2084[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2085 = {1{`RANDOM}};
  _T_6887_2022 = _RAND_2085[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2086 = {1{`RANDOM}};
  _T_6887_2023 = _RAND_2086[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2087 = {1{`RANDOM}};
  _T_6887_2024 = _RAND_2087[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2088 = {1{`RANDOM}};
  _T_6887_2025 = _RAND_2088[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2089 = {1{`RANDOM}};
  _T_6887_2026 = _RAND_2089[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2090 = {1{`RANDOM}};
  _T_6887_2027 = _RAND_2090[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2091 = {1{`RANDOM}};
  _T_6887_2028 = _RAND_2091[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2092 = {1{`RANDOM}};
  _T_6887_2029 = _RAND_2092[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2093 = {1{`RANDOM}};
  _T_6887_2030 = _RAND_2093[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2094 = {1{`RANDOM}};
  _T_6887_2031 = _RAND_2094[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2095 = {1{`RANDOM}};
  _T_6887_2032 = _RAND_2095[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2096 = {1{`RANDOM}};
  _T_6887_2033 = _RAND_2096[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2097 = {1{`RANDOM}};
  _T_6887_2034 = _RAND_2097[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2098 = {1{`RANDOM}};
  _T_6887_2035 = _RAND_2098[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2099 = {1{`RANDOM}};
  _T_6887_2036 = _RAND_2099[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2100 = {1{`RANDOM}};
  _T_6887_2037 = _RAND_2100[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2101 = {1{`RANDOM}};
  _T_6887_2038 = _RAND_2101[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2102 = {1{`RANDOM}};
  _T_6887_2039 = _RAND_2102[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2103 = {1{`RANDOM}};
  _T_6887_2040 = _RAND_2103[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2104 = {1{`RANDOM}};
  _T_6887_2041 = _RAND_2104[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2105 = {1{`RANDOM}};
  _T_6887_2042 = _RAND_2105[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2106 = {1{`RANDOM}};
  _T_6887_2043 = _RAND_2106[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2107 = {1{`RANDOM}};
  _T_6887_2044 = _RAND_2107[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2108 = {1{`RANDOM}};
  _T_6887_2045 = _RAND_2108[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2109 = {1{`RANDOM}};
  _T_6887_2046 = _RAND_2109[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2110 = {1{`RANDOM}};
  _T_6887_2047 = _RAND_2110[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2111 = {1{`RANDOM}};
  _T_13304_0 = _RAND_2111[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2112 = {1{`RANDOM}};
  _T_13304_1 = _RAND_2112[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2113 = {1{`RANDOM}};
  _T_13304_2 = _RAND_2113[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2114 = {1{`RANDOM}};
  _T_13304_3 = _RAND_2114[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2115 = {1{`RANDOM}};
  _T_13304_4 = _RAND_2115[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2116 = {1{`RANDOM}};
  _T_13304_5 = _RAND_2116[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2117 = {1{`RANDOM}};
  _T_13304_6 = _RAND_2117[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2118 = {1{`RANDOM}};
  _T_13304_7 = _RAND_2118[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2119 = {1{`RANDOM}};
  _T_13304_8 = _RAND_2119[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2120 = {1{`RANDOM}};
  _T_13304_9 = _RAND_2120[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2121 = {1{`RANDOM}};
  _T_13304_10 = _RAND_2121[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2122 = {1{`RANDOM}};
  _T_13304_11 = _RAND_2122[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2123 = {1{`RANDOM}};
  _T_13304_12 = _RAND_2123[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2124 = {1{`RANDOM}};
  _T_13304_13 = _RAND_2124[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2125 = {1{`RANDOM}};
  _T_13304_14 = _RAND_2125[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2126 = {1{`RANDOM}};
  _T_13304_15 = _RAND_2126[14:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2127 = {1{`RANDOM}};
  _T_13893 = _RAND_2127[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2128 = {1{`RANDOM}};
  value_1 = _RAND_2128[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2129 = {2{`RANDOM}};
  _T_14075_7 = _RAND_2129[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2130 = {2{`RANDOM}};
  _T_14075_6 = _RAND_2130[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2131 = {2{`RANDOM}};
  _T_14075_5 = _RAND_2131[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2132 = {2{`RANDOM}};
  _T_14075_4 = _RAND_2132[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2133 = {2{`RANDOM}};
  _T_14075_3 = _RAND_2133[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2134 = {2{`RANDOM}};
  _T_14075_2 = _RAND_2134[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2135 = {2{`RANDOM}};
  _T_14075_1 = _RAND_2135[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2136 = {2{`RANDOM}};
  _T_14075_0 = _RAND_2136[63:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2137 = {1{`RANDOM}};
  value_2 = _RAND_2137[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2138 = {1{`RANDOM}};
  value_3 = _RAND_2138[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      _T_258 <= 13'h0;
    end else begin
      if (_T_262) begin
        _T_258 <= _T_264;
      end
    end
    if (reset) begin
      _T_267 <= 4'h0;
    end else begin
      if (_T_14272) begin
        if (_T_321) begin
          _T_267 <= 4'h0;
        end else begin
          if (_T_14197) begin
            if (_T_14195) begin
              if (_T_301) begin
                _T_267 <= 4'h9;
              end else begin
                _T_267 <= 4'h7;
              end
            end else begin
              if (_T_14188) begin
                _T_267 <= 4'he;
              end else begin
                if (_T_14182) begin
                  if (_T_14098) begin
                    _T_267 <= 4'hd;
                  end else begin
                    if (_T_14179) begin
                      _T_267 <= 4'hc;
                    end else begin
                      if (_T_14170) begin
                        _T_267 <= 4'hb;
                      end else begin
                        if (_T_14162) begin
                          if (_T_301) begin
                            _T_267 <= 4'hf;
                          end else begin
                            _T_267 <= 4'h0;
                          end
                        end else begin
                          if (_T_14102) begin
                            if (_T_318) begin
                              _T_267 <= 4'h9;
                            end else begin
                              if (_T_13896) begin
                                if (_T_14097) begin
                                  if (_T_13153) begin
                                    _T_267 <= 4'hf;
                                  end else begin
                                    if (_T_14098) begin
                                      _T_267 <= 4'ha;
                                    end else begin
                                      if (_T_13154) begin
                                        _T_267 <= 4'h7;
                                      end else begin
                                        if (_T_482) begin
                                          if (_T_13383) begin
                                            _T_267 <= 4'h8;
                                          end else begin
                                            if (_T_13392) begin
                                              _T_267 <= 4'hd;
                                            end else begin
                                              if (_T_13036) begin
                                                _T_267 <= 4'h6;
                                              end else begin
                                                if (_T_484) begin
                                                  _T_267 <= 4'h5;
                                                end else begin
                                                  if (_T_458) begin
                                                    _T_267 <= 4'h4;
                                                  end else begin
                                                    if (_T_429) begin
                                                      if (_T_315) begin
                                                        _T_267 <= 4'h2;
                                                      end else begin
                                                        if (_T_335) begin
                                                          if (_T_284) begin
                                                            _T_267 <= 4'h4;
                                                          end else begin
                                                            if (_T_288) begin
                                                              _T_267 <= 4'h1;
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end else begin
                                                      if (_T_335) begin
                                                        if (_T_284) begin
                                                          _T_267 <= 4'h4;
                                                        end else begin
                                                          if (_T_288) begin
                                                            _T_267 <= 4'h1;
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end else begin
                                          if (_T_13036) begin
                                            _T_267 <= 4'h6;
                                          end else begin
                                            if (_T_484) begin
                                              _T_267 <= 4'h5;
                                            end else begin
                                              if (_T_458) begin
                                                _T_267 <= 4'h4;
                                              end else begin
                                                if (_T_429) begin
                                                  if (_T_315) begin
                                                    _T_267 <= 4'h2;
                                                  end else begin
                                                    if (_T_335) begin
                                                      if (_T_284) begin
                                                        _T_267 <= 4'h4;
                                                      end else begin
                                                        if (_T_288) begin
                                                          _T_267 <= 4'h1;
                                                        end
                                                      end
                                                    end
                                                  end
                                                end else begin
                                                  if (_T_335) begin
                                                    if (_T_284) begin
                                                      _T_267 <= 4'h4;
                                                    end else begin
                                                      if (_T_288) begin
                                                        _T_267 <= 4'h1;
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end else begin
                                  if (_T_482) begin
                                    if (_T_13383) begin
                                      _T_267 <= 4'h8;
                                    end else begin
                                      if (_T_13392) begin
                                        _T_267 <= 4'hd;
                                      end else begin
                                        if (_T_13036) begin
                                          _T_267 <= 4'h6;
                                        end else begin
                                          if (_T_484) begin
                                            _T_267 <= 4'h5;
                                          end else begin
                                            if (_T_458) begin
                                              _T_267 <= 4'h4;
                                            end else begin
                                              if (_T_429) begin
                                                if (_T_315) begin
                                                  _T_267 <= 4'h2;
                                                end else begin
                                                  _T_267 <= _GEN_35;
                                                end
                                              end else begin
                                                _T_267 <= _GEN_35;
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end else begin
                                    if (_T_13036) begin
                                      _T_267 <= 4'h6;
                                    end else begin
                                      if (_T_484) begin
                                        _T_267 <= 4'h5;
                                      end else begin
                                        if (_T_458) begin
                                          _T_267 <= 4'h4;
                                        end else begin
                                          if (_T_429) begin
                                            if (_T_315) begin
                                              _T_267 <= 4'h2;
                                            end else begin
                                              _T_267 <= _GEN_35;
                                            end
                                          end else begin
                                            _T_267 <= _GEN_35;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end else begin
                                if (_T_482) begin
                                  if (_T_13383) begin
                                    _T_267 <= 4'h8;
                                  end else begin
                                    if (_T_13392) begin
                                      _T_267 <= 4'hd;
                                    end else begin
                                      _T_267 <= _GEN_4175;
                                    end
                                  end
                                end else begin
                                  _T_267 <= _GEN_4175;
                                end
                              end
                            end
                          end else begin
                            if (_T_13896) begin
                              if (_T_14097) begin
                                if (_T_13153) begin
                                  _T_267 <= 4'hf;
                                end else begin
                                  if (_T_14098) begin
                                    _T_267 <= 4'ha;
                                  end else begin
                                    if (_T_13154) begin
                                      _T_267 <= 4'h7;
                                    end else begin
                                      if (_T_482) begin
                                        if (_T_13383) begin
                                          _T_267 <= 4'h8;
                                        end else begin
                                          if (_T_13392) begin
                                            _T_267 <= 4'hd;
                                          end else begin
                                            _T_267 <= _GEN_4175;
                                          end
                                        end
                                      end else begin
                                        _T_267 <= _GEN_4175;
                                      end
                                    end
                                  end
                                end
                              end else begin
                                _T_267 <= _GEN_6309;
                              end
                            end else begin
                              _T_267 <= _GEN_6309;
                            end
                          end
                        end
                      end
                    end
                  end
                end else begin
                  if (_T_14179) begin
                    _T_267 <= 4'hc;
                  end else begin
                    if (_T_14170) begin
                      _T_267 <= 4'hb;
                    end else begin
                      if (_T_14162) begin
                        if (_T_301) begin
                          _T_267 <= 4'hf;
                        end else begin
                          _T_267 <= 4'h0;
                        end
                      end else begin
                        if (_T_14102) begin
                          if (_T_318) begin
                            _T_267 <= 4'h9;
                          end else begin
                            if (_T_13896) begin
                              if (_T_14097) begin
                                if (_T_13153) begin
                                  _T_267 <= 4'hf;
                                end else begin
                                  if (_T_14098) begin
                                    _T_267 <= 4'ha;
                                  end else begin
                                    if (_T_13154) begin
                                      _T_267 <= 4'h7;
                                    end else begin
                                      _T_267 <= _GEN_6309;
                                    end
                                  end
                                end
                              end else begin
                                _T_267 <= _GEN_6309;
                              end
                            end else begin
                              _T_267 <= _GEN_6309;
                            end
                          end
                        end else begin
                          if (_T_13896) begin
                            if (_T_14097) begin
                              if (_T_13153) begin
                                _T_267 <= 4'hf;
                              end else begin
                                if (_T_14098) begin
                                  _T_267 <= 4'ha;
                                end else begin
                                  if (_T_13154) begin
                                    _T_267 <= 4'h7;
                                  end else begin
                                    _T_267 <= _GEN_6309;
                                  end
                                end
                              end
                            end else begin
                              _T_267 <= _GEN_6309;
                            end
                          end else begin
                            _T_267 <= _GEN_6309;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end else begin
            if (_T_14188) begin
              _T_267 <= 4'he;
            end else begin
              if (_T_14182) begin
                if (_T_14098) begin
                  _T_267 <= 4'hd;
                end else begin
                  if (_T_14179) begin
                    _T_267 <= 4'hc;
                  end else begin
                    if (_T_14170) begin
                      _T_267 <= 4'hb;
                    end else begin
                      if (_T_14162) begin
                        if (_T_301) begin
                          _T_267 <= 4'hf;
                        end else begin
                          _T_267 <= 4'h0;
                        end
                      end else begin
                        if (_T_14102) begin
                          if (_T_318) begin
                            _T_267 <= 4'h9;
                          end else begin
                            _T_267 <= _GEN_6922;
                          end
                        end else begin
                          _T_267 <= _GEN_6922;
                        end
                      end
                    end
                  end
                end
              end else begin
                if (_T_14179) begin
                  _T_267 <= 4'hc;
                end else begin
                  if (_T_14170) begin
                    _T_267 <= 4'hb;
                  end else begin
                    if (_T_14162) begin
                      if (_T_301) begin
                        _T_267 <= 4'hf;
                      end else begin
                        _T_267 <= 4'h0;
                      end
                    end else begin
                      if (_T_14102) begin
                        if (_T_318) begin
                          _T_267 <= 4'h9;
                        end else begin
                          _T_267 <= _GEN_6922;
                        end
                      end else begin
                        _T_267 <= _GEN_6922;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_14197) begin
          if (_T_14195) begin
            if (_T_301) begin
              _T_267 <= 4'h9;
            end else begin
              _T_267 <= 4'h7;
            end
          end else begin
            if (_T_14188) begin
              _T_267 <= 4'he;
            end else begin
              if (_T_14182) begin
                if (_T_14098) begin
                  _T_267 <= 4'hd;
                end else begin
                  _T_267 <= _GEN_6979;
                end
              end else begin
                _T_267 <= _GEN_6979;
              end
            end
          end
        end else begin
          if (_T_14188) begin
            _T_267 <= 4'he;
          end else begin
            if (_T_14182) begin
              if (_T_14098) begin
                _T_267 <= 4'hd;
              end else begin
                _T_267 <= _GEN_6979;
              end
            end else begin
              _T_267 <= _GEN_6979;
            end
          end
        end
      end
    end
    if (_T_335) begin
      if (_T_284) begin
        _T_291 <= auto_in_a_bits_address;
      end else begin
        if (_T_288) begin
          _T_291 <= auto_in_a_bits_address;
        end
      end
    end
    if (_T_335) begin
      if (_T_284) begin
        _T_293 <= auto_in_a_bits_source;
      end else begin
        if (_T_288) begin
          _T_293 <= auto_in_a_bits_source;
        end
      end
    end
    if (reset) begin
      _T_297 <= 4'hf;
    end else begin
      _T_297 <= _GEN_30[3:0];
    end
    if (_T_335) begin
      if (_T_284) begin
        _T_299 <= auto_in_a_bits_size;
      end else begin
        if (_T_288) begin
          _T_299 <= auto_in_a_bits_size;
        end
      end
    end
    if (reset) begin
      _T_301 <= 1'h0;
    end else begin
      if (_T_335) begin
        if (_T_284) begin
          _T_301 <= 1'h1;
        end else begin
          if (_T_288) begin
            _T_301 <= 1'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_303 <= 1'h0;
    end else begin
      if (_T_335) begin
        if (_T_284) begin
          _T_303 <= 1'h0;
        end else begin
          if (_T_288) begin
            _T_303 <= 1'h1;
          end
        end
      end
    end
    _T_306 <= _GEN_34[3:0];
    if (reset) begin
      _T_312 <= 3'h0;
    end else begin
      if (_T_429) begin
        if (_T_335) begin
          _T_312 <= _T_432;
        end else begin
          if (_T_426) begin
            _T_312 <= _T_435;
          end
        end
      end
    end
    if (reset) begin
      _T_317 <= 3'h0;
    end else begin
      if (_T_14102) begin
        _T_317 <= _T_14104;
      end else begin
        if (_T_335) begin
          if (_T_284) begin
            _T_317 <= _T_304;
          end else begin
            if (_T_288) begin
              _T_317 <= _T_304;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_320 <= 3'h0;
    end else begin
      if (_T_14272) begin
        _T_320 <= _T_14274;
      end else begin
        if (_T_335) begin
          if (_T_284) begin
            _T_320 <= _T_304;
          end else begin
            if (_T_288) begin
              _T_320 <= _T_304;
            end
          end
        end
      end
    end
    if (_T_429) begin
      if (3'h0 == _T_441) begin
        _T_344_0 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h1 == _T_441) begin
        _T_344_1 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h2 == _T_441) begin
        _T_344_2 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h3 == _T_441) begin
        _T_344_3 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h4 == _T_441) begin
        _T_344_4 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h5 == _T_441) begin
        _T_344_5 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h6 == _T_441) begin
        _T_344_6 <= auto_in_a_bits_data;
      end
    end
    if (_T_429) begin
      if (3'h7 == _T_441) begin
        _T_344_7 <= auto_in_a_bits_data;
      end
    end
    if (reset) begin
      _T_397_0 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h0 == _T_441) begin
          _T_397_0 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_1 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h1 == _T_441) begin
          _T_397_1 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_2 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h2 == _T_441) begin
          _T_397_2 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_3 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h3 == _T_441) begin
          _T_397_3 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_4 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h4 == _T_441) begin
          _T_397_4 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_5 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h5 == _T_441) begin
          _T_397_5 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_6 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h6 == _T_441) begin
          _T_397_6 <= auto_in_a_bits_mask;
        end
      end
    end
    if (reset) begin
      _T_397_7 <= 8'h0;
    end else begin
      if (_T_429) begin
        if (3'h7 == _T_441) begin
          _T_397_7 <= auto_in_a_bits_mask;
        end
      end
    end
    if (_T_13036) begin
      _T_684 <= _T_563;
    end
    if (_T_13036) begin
      _T_686 <= _T_600;
    end
    if (_T_13036) begin
      _T_690_0 <= _T_604_0;
    end
    if (_T_13036) begin
      _T_690_1 <= _T_604_1;
    end
    if (_T_13036) begin
      _T_690_2 <= _T_604_2;
    end
    if (_T_13036) begin
      _T_690_3 <= _T_604_3;
    end
    if (_T_13036) begin
      _T_690_4 <= _T_604_4;
    end
    if (_T_13036) begin
      _T_690_5 <= _T_604_5;
    end
    if (_T_13036) begin
      _T_690_6 <= _T_604_6;
    end
    if (_T_13036) begin
      _T_690_7 <= _T_604_7;
    end
    if (_T_13036) begin
      _T_690_8 <= _T_604_8;
    end
    if (_T_13036) begin
      _T_690_9 <= _T_604_9;
    end
    if (_T_13036) begin
      _T_690_10 <= _T_604_10;
    end
    if (_T_13036) begin
      _T_690_11 <= _T_604_11;
    end
    if (_T_13036) begin
      _T_690_12 <= _T_604_12;
    end
    if (_T_13036) begin
      _T_690_13 <= _T_604_13;
    end
    if (_T_13036) begin
      _T_690_14 <= _T_604_14;
    end
    if (_T_13036) begin
      _T_690_15 <= _T_604_15;
    end
    if (_T_13036) begin
      if (_GEN_2126) begin
        _T_710 <= 16'hffff;
      end else begin
        _T_710 <= _T_659;
      end
    end
    if (_T_13036) begin
      _T_714_0 <= _T_663_0;
    end
    if (_T_13036) begin
      _T_714_1 <= _T_663_1;
    end
    if (_T_13036) begin
      _T_714_2 <= _T_663_2;
    end
    if (_T_13036) begin
      _T_714_3 <= _T_663_3;
    end
    if (_T_13036) begin
      _T_714_4 <= _T_663_4;
    end
    if (_T_13036) begin
      _T_714_5 <= _T_663_5;
    end
    if (_T_13036) begin
      _T_714_6 <= _T_663_6;
    end
    if (_T_13036) begin
      _T_714_7 <= _T_663_7;
    end
    if (_T_13036) begin
      _T_714_8 <= _T_663_8;
    end
    if (_T_13036) begin
      _T_714_9 <= _T_663_9;
    end
    if (_T_13036) begin
      _T_714_10 <= _T_663_10;
    end
    if (_T_13036) begin
      _T_714_11 <= _T_663_11;
    end
    if (_T_13036) begin
      _T_714_12 <= _T_663_12;
    end
    if (_T_13036) begin
      _T_714_13 <= _T_663_13;
    end
    if (_T_13036) begin
      _T_714_14 <= _T_663_14;
    end
    if (_T_13036) begin
      _T_714_15 <= _T_663_15;
    end
    if (reset) begin
      _T_6887_0 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h0 == _T_481) begin
          _T_6887_0 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1 == _T_481) begin
          _T_6887_1 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2 == _T_481) begin
          _T_6887_2 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_3 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3 == _T_481) begin
          _T_6887_3 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_4 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4 == _T_481) begin
          _T_6887_4 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_5 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5 == _T_481) begin
          _T_6887_5 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_6 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6 == _T_481) begin
          _T_6887_6 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_7 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7 == _T_481) begin
          _T_6887_7 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_8 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8 == _T_481) begin
          _T_6887_8 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_9 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9 == _T_481) begin
          _T_6887_9 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_10 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha == _T_481) begin
          _T_6887_10 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_11 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb == _T_481) begin
          _T_6887_11 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_12 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc == _T_481) begin
          _T_6887_12 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_13 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd == _T_481) begin
          _T_6887_13 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_14 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he == _T_481) begin
          _T_6887_14 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_15 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf == _T_481) begin
          _T_6887_15 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_16 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10 == _T_481) begin
          _T_6887_16 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_17 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11 == _T_481) begin
          _T_6887_17 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_18 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12 == _T_481) begin
          _T_6887_18 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_19 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13 == _T_481) begin
          _T_6887_19 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_20 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14 == _T_481) begin
          _T_6887_20 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_21 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15 == _T_481) begin
          _T_6887_21 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_22 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16 == _T_481) begin
          _T_6887_22 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_23 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17 == _T_481) begin
          _T_6887_23 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_24 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18 == _T_481) begin
          _T_6887_24 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_25 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19 == _T_481) begin
          _T_6887_25 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_26 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a == _T_481) begin
          _T_6887_26 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_27 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b == _T_481) begin
          _T_6887_27 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_28 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c == _T_481) begin
          _T_6887_28 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_29 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d == _T_481) begin
          _T_6887_29 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_30 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e == _T_481) begin
          _T_6887_30 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_31 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f == _T_481) begin
          _T_6887_31 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_32 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20 == _T_481) begin
          _T_6887_32 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_33 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21 == _T_481) begin
          _T_6887_33 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_34 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22 == _T_481) begin
          _T_6887_34 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_35 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23 == _T_481) begin
          _T_6887_35 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_36 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24 == _T_481) begin
          _T_6887_36 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_37 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25 == _T_481) begin
          _T_6887_37 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_38 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26 == _T_481) begin
          _T_6887_38 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_39 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27 == _T_481) begin
          _T_6887_39 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_40 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28 == _T_481) begin
          _T_6887_40 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_41 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29 == _T_481) begin
          _T_6887_41 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_42 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a == _T_481) begin
          _T_6887_42 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_43 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b == _T_481) begin
          _T_6887_43 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_44 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c == _T_481) begin
          _T_6887_44 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_45 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d == _T_481) begin
          _T_6887_45 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_46 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e == _T_481) begin
          _T_6887_46 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_47 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f == _T_481) begin
          _T_6887_47 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_48 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30 == _T_481) begin
          _T_6887_48 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_49 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31 == _T_481) begin
          _T_6887_49 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_50 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32 == _T_481) begin
          _T_6887_50 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_51 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33 == _T_481) begin
          _T_6887_51 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_52 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34 == _T_481) begin
          _T_6887_52 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_53 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35 == _T_481) begin
          _T_6887_53 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_54 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36 == _T_481) begin
          _T_6887_54 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_55 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37 == _T_481) begin
          _T_6887_55 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_56 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38 == _T_481) begin
          _T_6887_56 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_57 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39 == _T_481) begin
          _T_6887_57 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_58 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a == _T_481) begin
          _T_6887_58 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_59 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b == _T_481) begin
          _T_6887_59 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_60 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c == _T_481) begin
          _T_6887_60 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_61 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d == _T_481) begin
          _T_6887_61 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_62 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e == _T_481) begin
          _T_6887_62 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_63 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f == _T_481) begin
          _T_6887_63 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_64 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40 == _T_481) begin
          _T_6887_64 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_65 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41 == _T_481) begin
          _T_6887_65 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_66 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42 == _T_481) begin
          _T_6887_66 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_67 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43 == _T_481) begin
          _T_6887_67 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_68 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44 == _T_481) begin
          _T_6887_68 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_69 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45 == _T_481) begin
          _T_6887_69 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_70 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46 == _T_481) begin
          _T_6887_70 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_71 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47 == _T_481) begin
          _T_6887_71 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_72 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48 == _T_481) begin
          _T_6887_72 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_73 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49 == _T_481) begin
          _T_6887_73 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_74 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a == _T_481) begin
          _T_6887_74 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_75 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b == _T_481) begin
          _T_6887_75 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_76 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c == _T_481) begin
          _T_6887_76 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_77 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d == _T_481) begin
          _T_6887_77 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_78 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e == _T_481) begin
          _T_6887_78 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_79 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f == _T_481) begin
          _T_6887_79 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_80 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50 == _T_481) begin
          _T_6887_80 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_81 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51 == _T_481) begin
          _T_6887_81 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_82 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52 == _T_481) begin
          _T_6887_82 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_83 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53 == _T_481) begin
          _T_6887_83 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_84 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54 == _T_481) begin
          _T_6887_84 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_85 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55 == _T_481) begin
          _T_6887_85 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_86 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56 == _T_481) begin
          _T_6887_86 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_87 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57 == _T_481) begin
          _T_6887_87 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_88 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58 == _T_481) begin
          _T_6887_88 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_89 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59 == _T_481) begin
          _T_6887_89 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_90 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a == _T_481) begin
          _T_6887_90 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_91 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b == _T_481) begin
          _T_6887_91 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_92 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c == _T_481) begin
          _T_6887_92 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_93 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d == _T_481) begin
          _T_6887_93 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_94 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e == _T_481) begin
          _T_6887_94 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_95 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f == _T_481) begin
          _T_6887_95 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_96 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60 == _T_481) begin
          _T_6887_96 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_97 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61 == _T_481) begin
          _T_6887_97 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_98 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62 == _T_481) begin
          _T_6887_98 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_99 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63 == _T_481) begin
          _T_6887_99 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_100 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64 == _T_481) begin
          _T_6887_100 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_101 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65 == _T_481) begin
          _T_6887_101 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_102 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66 == _T_481) begin
          _T_6887_102 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_103 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67 == _T_481) begin
          _T_6887_103 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_104 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68 == _T_481) begin
          _T_6887_104 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_105 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69 == _T_481) begin
          _T_6887_105 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_106 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a == _T_481) begin
          _T_6887_106 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_107 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b == _T_481) begin
          _T_6887_107 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_108 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c == _T_481) begin
          _T_6887_108 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_109 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d == _T_481) begin
          _T_6887_109 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_110 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e == _T_481) begin
          _T_6887_110 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_111 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f == _T_481) begin
          _T_6887_111 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_112 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70 == _T_481) begin
          _T_6887_112 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_113 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71 == _T_481) begin
          _T_6887_113 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_114 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72 == _T_481) begin
          _T_6887_114 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_115 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73 == _T_481) begin
          _T_6887_115 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_116 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74 == _T_481) begin
          _T_6887_116 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_117 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75 == _T_481) begin
          _T_6887_117 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_118 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76 == _T_481) begin
          _T_6887_118 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_119 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77 == _T_481) begin
          _T_6887_119 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_120 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78 == _T_481) begin
          _T_6887_120 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_121 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79 == _T_481) begin
          _T_6887_121 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_122 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a == _T_481) begin
          _T_6887_122 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_123 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b == _T_481) begin
          _T_6887_123 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_124 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c == _T_481) begin
          _T_6887_124 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_125 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d == _T_481) begin
          _T_6887_125 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_126 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e == _T_481) begin
          _T_6887_126 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_127 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f == _T_481) begin
          _T_6887_127 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_128 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h80 == _T_481) begin
          _T_6887_128 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_129 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h81 == _T_481) begin
          _T_6887_129 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_130 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h82 == _T_481) begin
          _T_6887_130 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_131 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h83 == _T_481) begin
          _T_6887_131 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_132 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h84 == _T_481) begin
          _T_6887_132 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_133 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h85 == _T_481) begin
          _T_6887_133 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_134 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h86 == _T_481) begin
          _T_6887_134 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_135 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h87 == _T_481) begin
          _T_6887_135 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_136 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h88 == _T_481) begin
          _T_6887_136 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_137 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h89 == _T_481) begin
          _T_6887_137 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_138 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8a == _T_481) begin
          _T_6887_138 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_139 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8b == _T_481) begin
          _T_6887_139 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_140 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8c == _T_481) begin
          _T_6887_140 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_141 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8d == _T_481) begin
          _T_6887_141 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_142 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8e == _T_481) begin
          _T_6887_142 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_143 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h8f == _T_481) begin
          _T_6887_143 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_144 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h90 == _T_481) begin
          _T_6887_144 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_145 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h91 == _T_481) begin
          _T_6887_145 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_146 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h92 == _T_481) begin
          _T_6887_146 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_147 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h93 == _T_481) begin
          _T_6887_147 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_148 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h94 == _T_481) begin
          _T_6887_148 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_149 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h95 == _T_481) begin
          _T_6887_149 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_150 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h96 == _T_481) begin
          _T_6887_150 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_151 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h97 == _T_481) begin
          _T_6887_151 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_152 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h98 == _T_481) begin
          _T_6887_152 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_153 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h99 == _T_481) begin
          _T_6887_153 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_154 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9a == _T_481) begin
          _T_6887_154 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_155 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9b == _T_481) begin
          _T_6887_155 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_156 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9c == _T_481) begin
          _T_6887_156 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_157 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9d == _T_481) begin
          _T_6887_157 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_158 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9e == _T_481) begin
          _T_6887_158 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_159 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h9f == _T_481) begin
          _T_6887_159 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_160 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha0 == _T_481) begin
          _T_6887_160 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_161 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha1 == _T_481) begin
          _T_6887_161 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_162 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha2 == _T_481) begin
          _T_6887_162 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_163 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha3 == _T_481) begin
          _T_6887_163 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_164 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha4 == _T_481) begin
          _T_6887_164 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_165 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha5 == _T_481) begin
          _T_6887_165 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_166 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha6 == _T_481) begin
          _T_6887_166 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_167 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha7 == _T_481) begin
          _T_6887_167 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_168 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha8 == _T_481) begin
          _T_6887_168 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_169 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'ha9 == _T_481) begin
          _T_6887_169 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_170 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'haa == _T_481) begin
          _T_6887_170 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_171 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hab == _T_481) begin
          _T_6887_171 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_172 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hac == _T_481) begin
          _T_6887_172 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_173 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'had == _T_481) begin
          _T_6887_173 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_174 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hae == _T_481) begin
          _T_6887_174 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_175 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'haf == _T_481) begin
          _T_6887_175 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_176 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb0 == _T_481) begin
          _T_6887_176 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_177 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb1 == _T_481) begin
          _T_6887_177 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_178 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb2 == _T_481) begin
          _T_6887_178 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_179 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb3 == _T_481) begin
          _T_6887_179 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_180 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb4 == _T_481) begin
          _T_6887_180 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_181 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb5 == _T_481) begin
          _T_6887_181 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_182 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb6 == _T_481) begin
          _T_6887_182 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_183 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb7 == _T_481) begin
          _T_6887_183 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_184 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb8 == _T_481) begin
          _T_6887_184 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_185 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hb9 == _T_481) begin
          _T_6887_185 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_186 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hba == _T_481) begin
          _T_6887_186 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_187 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hbb == _T_481) begin
          _T_6887_187 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_188 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hbc == _T_481) begin
          _T_6887_188 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_189 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hbd == _T_481) begin
          _T_6887_189 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_190 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hbe == _T_481) begin
          _T_6887_190 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_191 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hbf == _T_481) begin
          _T_6887_191 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_192 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc0 == _T_481) begin
          _T_6887_192 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_193 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc1 == _T_481) begin
          _T_6887_193 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_194 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc2 == _T_481) begin
          _T_6887_194 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_195 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc3 == _T_481) begin
          _T_6887_195 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_196 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc4 == _T_481) begin
          _T_6887_196 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_197 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc5 == _T_481) begin
          _T_6887_197 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_198 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc6 == _T_481) begin
          _T_6887_198 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_199 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc7 == _T_481) begin
          _T_6887_199 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_200 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc8 == _T_481) begin
          _T_6887_200 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_201 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hc9 == _T_481) begin
          _T_6887_201 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_202 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hca == _T_481) begin
          _T_6887_202 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_203 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hcb == _T_481) begin
          _T_6887_203 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_204 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hcc == _T_481) begin
          _T_6887_204 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_205 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hcd == _T_481) begin
          _T_6887_205 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_206 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hce == _T_481) begin
          _T_6887_206 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_207 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hcf == _T_481) begin
          _T_6887_207 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_208 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd0 == _T_481) begin
          _T_6887_208 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_209 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd1 == _T_481) begin
          _T_6887_209 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_210 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd2 == _T_481) begin
          _T_6887_210 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_211 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd3 == _T_481) begin
          _T_6887_211 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_212 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd4 == _T_481) begin
          _T_6887_212 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_213 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd5 == _T_481) begin
          _T_6887_213 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_214 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd6 == _T_481) begin
          _T_6887_214 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_215 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd7 == _T_481) begin
          _T_6887_215 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_216 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd8 == _T_481) begin
          _T_6887_216 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_217 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hd9 == _T_481) begin
          _T_6887_217 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_218 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hda == _T_481) begin
          _T_6887_218 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_219 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hdb == _T_481) begin
          _T_6887_219 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_220 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hdc == _T_481) begin
          _T_6887_220 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_221 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hdd == _T_481) begin
          _T_6887_221 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_222 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hde == _T_481) begin
          _T_6887_222 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_223 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hdf == _T_481) begin
          _T_6887_223 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_224 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he0 == _T_481) begin
          _T_6887_224 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_225 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he1 == _T_481) begin
          _T_6887_225 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_226 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he2 == _T_481) begin
          _T_6887_226 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_227 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he3 == _T_481) begin
          _T_6887_227 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_228 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he4 == _T_481) begin
          _T_6887_228 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_229 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he5 == _T_481) begin
          _T_6887_229 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_230 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he6 == _T_481) begin
          _T_6887_230 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_231 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he7 == _T_481) begin
          _T_6887_231 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_232 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he8 == _T_481) begin
          _T_6887_232 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_233 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'he9 == _T_481) begin
          _T_6887_233 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_234 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hea == _T_481) begin
          _T_6887_234 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_235 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'heb == _T_481) begin
          _T_6887_235 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_236 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hec == _T_481) begin
          _T_6887_236 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_237 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hed == _T_481) begin
          _T_6887_237 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_238 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hee == _T_481) begin
          _T_6887_238 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_239 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hef == _T_481) begin
          _T_6887_239 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_240 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf0 == _T_481) begin
          _T_6887_240 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_241 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf1 == _T_481) begin
          _T_6887_241 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_242 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf2 == _T_481) begin
          _T_6887_242 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_243 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf3 == _T_481) begin
          _T_6887_243 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_244 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf4 == _T_481) begin
          _T_6887_244 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_245 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf5 == _T_481) begin
          _T_6887_245 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_246 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf6 == _T_481) begin
          _T_6887_246 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_247 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf7 == _T_481) begin
          _T_6887_247 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_248 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf8 == _T_481) begin
          _T_6887_248 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_249 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hf9 == _T_481) begin
          _T_6887_249 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_250 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hfa == _T_481) begin
          _T_6887_250 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_251 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hfb == _T_481) begin
          _T_6887_251 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_252 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hfc == _T_481) begin
          _T_6887_252 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_253 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hfd == _T_481) begin
          _T_6887_253 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_254 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hfe == _T_481) begin
          _T_6887_254 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_255 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'hff == _T_481) begin
          _T_6887_255 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_256 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h100 == _T_481) begin
          _T_6887_256 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_257 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h101 == _T_481) begin
          _T_6887_257 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_258 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h102 == _T_481) begin
          _T_6887_258 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_259 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h103 == _T_481) begin
          _T_6887_259 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_260 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h104 == _T_481) begin
          _T_6887_260 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_261 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h105 == _T_481) begin
          _T_6887_261 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_262 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h106 == _T_481) begin
          _T_6887_262 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_263 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h107 == _T_481) begin
          _T_6887_263 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_264 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h108 == _T_481) begin
          _T_6887_264 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_265 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h109 == _T_481) begin
          _T_6887_265 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_266 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10a == _T_481) begin
          _T_6887_266 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_267 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10b == _T_481) begin
          _T_6887_267 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_268 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10c == _T_481) begin
          _T_6887_268 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_269 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10d == _T_481) begin
          _T_6887_269 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_270 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10e == _T_481) begin
          _T_6887_270 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_271 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h10f == _T_481) begin
          _T_6887_271 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_272 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h110 == _T_481) begin
          _T_6887_272 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_273 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h111 == _T_481) begin
          _T_6887_273 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_274 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h112 == _T_481) begin
          _T_6887_274 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_275 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h113 == _T_481) begin
          _T_6887_275 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_276 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h114 == _T_481) begin
          _T_6887_276 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_277 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h115 == _T_481) begin
          _T_6887_277 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_278 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h116 == _T_481) begin
          _T_6887_278 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_279 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h117 == _T_481) begin
          _T_6887_279 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_280 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h118 == _T_481) begin
          _T_6887_280 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_281 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h119 == _T_481) begin
          _T_6887_281 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_282 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11a == _T_481) begin
          _T_6887_282 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_283 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11b == _T_481) begin
          _T_6887_283 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_284 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11c == _T_481) begin
          _T_6887_284 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_285 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11d == _T_481) begin
          _T_6887_285 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_286 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11e == _T_481) begin
          _T_6887_286 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_287 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h11f == _T_481) begin
          _T_6887_287 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_288 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h120 == _T_481) begin
          _T_6887_288 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_289 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h121 == _T_481) begin
          _T_6887_289 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_290 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h122 == _T_481) begin
          _T_6887_290 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_291 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h123 == _T_481) begin
          _T_6887_291 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_292 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h124 == _T_481) begin
          _T_6887_292 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_293 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h125 == _T_481) begin
          _T_6887_293 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_294 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h126 == _T_481) begin
          _T_6887_294 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_295 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h127 == _T_481) begin
          _T_6887_295 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_296 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h128 == _T_481) begin
          _T_6887_296 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_297 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h129 == _T_481) begin
          _T_6887_297 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_298 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12a == _T_481) begin
          _T_6887_298 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_299 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12b == _T_481) begin
          _T_6887_299 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_300 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12c == _T_481) begin
          _T_6887_300 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_301 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12d == _T_481) begin
          _T_6887_301 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_302 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12e == _T_481) begin
          _T_6887_302 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_303 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h12f == _T_481) begin
          _T_6887_303 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_304 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h130 == _T_481) begin
          _T_6887_304 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_305 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h131 == _T_481) begin
          _T_6887_305 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_306 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h132 == _T_481) begin
          _T_6887_306 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_307 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h133 == _T_481) begin
          _T_6887_307 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_308 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h134 == _T_481) begin
          _T_6887_308 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_309 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h135 == _T_481) begin
          _T_6887_309 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_310 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h136 == _T_481) begin
          _T_6887_310 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_311 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h137 == _T_481) begin
          _T_6887_311 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_312 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h138 == _T_481) begin
          _T_6887_312 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_313 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h139 == _T_481) begin
          _T_6887_313 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_314 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13a == _T_481) begin
          _T_6887_314 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_315 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13b == _T_481) begin
          _T_6887_315 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_316 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13c == _T_481) begin
          _T_6887_316 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_317 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13d == _T_481) begin
          _T_6887_317 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_318 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13e == _T_481) begin
          _T_6887_318 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_319 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h13f == _T_481) begin
          _T_6887_319 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_320 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h140 == _T_481) begin
          _T_6887_320 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_321 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h141 == _T_481) begin
          _T_6887_321 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_322 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h142 == _T_481) begin
          _T_6887_322 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_323 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h143 == _T_481) begin
          _T_6887_323 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_324 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h144 == _T_481) begin
          _T_6887_324 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_325 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h145 == _T_481) begin
          _T_6887_325 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_326 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h146 == _T_481) begin
          _T_6887_326 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_327 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h147 == _T_481) begin
          _T_6887_327 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_328 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h148 == _T_481) begin
          _T_6887_328 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_329 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h149 == _T_481) begin
          _T_6887_329 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_330 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14a == _T_481) begin
          _T_6887_330 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_331 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14b == _T_481) begin
          _T_6887_331 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_332 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14c == _T_481) begin
          _T_6887_332 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_333 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14d == _T_481) begin
          _T_6887_333 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_334 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14e == _T_481) begin
          _T_6887_334 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_335 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h14f == _T_481) begin
          _T_6887_335 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_336 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h150 == _T_481) begin
          _T_6887_336 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_337 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h151 == _T_481) begin
          _T_6887_337 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_338 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h152 == _T_481) begin
          _T_6887_338 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_339 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h153 == _T_481) begin
          _T_6887_339 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_340 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h154 == _T_481) begin
          _T_6887_340 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_341 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h155 == _T_481) begin
          _T_6887_341 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_342 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h156 == _T_481) begin
          _T_6887_342 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_343 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h157 == _T_481) begin
          _T_6887_343 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_344 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h158 == _T_481) begin
          _T_6887_344 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_345 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h159 == _T_481) begin
          _T_6887_345 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_346 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15a == _T_481) begin
          _T_6887_346 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_347 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15b == _T_481) begin
          _T_6887_347 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_348 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15c == _T_481) begin
          _T_6887_348 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_349 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15d == _T_481) begin
          _T_6887_349 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_350 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15e == _T_481) begin
          _T_6887_350 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_351 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h15f == _T_481) begin
          _T_6887_351 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_352 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h160 == _T_481) begin
          _T_6887_352 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_353 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h161 == _T_481) begin
          _T_6887_353 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_354 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h162 == _T_481) begin
          _T_6887_354 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_355 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h163 == _T_481) begin
          _T_6887_355 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_356 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h164 == _T_481) begin
          _T_6887_356 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_357 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h165 == _T_481) begin
          _T_6887_357 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_358 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h166 == _T_481) begin
          _T_6887_358 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_359 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h167 == _T_481) begin
          _T_6887_359 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_360 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h168 == _T_481) begin
          _T_6887_360 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_361 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h169 == _T_481) begin
          _T_6887_361 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_362 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16a == _T_481) begin
          _T_6887_362 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_363 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16b == _T_481) begin
          _T_6887_363 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_364 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16c == _T_481) begin
          _T_6887_364 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_365 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16d == _T_481) begin
          _T_6887_365 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_366 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16e == _T_481) begin
          _T_6887_366 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_367 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h16f == _T_481) begin
          _T_6887_367 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_368 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h170 == _T_481) begin
          _T_6887_368 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_369 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h171 == _T_481) begin
          _T_6887_369 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_370 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h172 == _T_481) begin
          _T_6887_370 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_371 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h173 == _T_481) begin
          _T_6887_371 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_372 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h174 == _T_481) begin
          _T_6887_372 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_373 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h175 == _T_481) begin
          _T_6887_373 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_374 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h176 == _T_481) begin
          _T_6887_374 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_375 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h177 == _T_481) begin
          _T_6887_375 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_376 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h178 == _T_481) begin
          _T_6887_376 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_377 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h179 == _T_481) begin
          _T_6887_377 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_378 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17a == _T_481) begin
          _T_6887_378 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_379 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17b == _T_481) begin
          _T_6887_379 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_380 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17c == _T_481) begin
          _T_6887_380 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_381 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17d == _T_481) begin
          _T_6887_381 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_382 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17e == _T_481) begin
          _T_6887_382 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_383 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h17f == _T_481) begin
          _T_6887_383 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_384 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h180 == _T_481) begin
          _T_6887_384 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_385 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h181 == _T_481) begin
          _T_6887_385 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_386 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h182 == _T_481) begin
          _T_6887_386 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_387 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h183 == _T_481) begin
          _T_6887_387 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_388 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h184 == _T_481) begin
          _T_6887_388 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_389 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h185 == _T_481) begin
          _T_6887_389 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_390 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h186 == _T_481) begin
          _T_6887_390 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_391 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h187 == _T_481) begin
          _T_6887_391 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_392 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h188 == _T_481) begin
          _T_6887_392 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_393 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h189 == _T_481) begin
          _T_6887_393 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_394 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18a == _T_481) begin
          _T_6887_394 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_395 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18b == _T_481) begin
          _T_6887_395 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_396 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18c == _T_481) begin
          _T_6887_396 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_397 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18d == _T_481) begin
          _T_6887_397 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_398 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18e == _T_481) begin
          _T_6887_398 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_399 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h18f == _T_481) begin
          _T_6887_399 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_400 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h190 == _T_481) begin
          _T_6887_400 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_401 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h191 == _T_481) begin
          _T_6887_401 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_402 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h192 == _T_481) begin
          _T_6887_402 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_403 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h193 == _T_481) begin
          _T_6887_403 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_404 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h194 == _T_481) begin
          _T_6887_404 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_405 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h195 == _T_481) begin
          _T_6887_405 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_406 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h196 == _T_481) begin
          _T_6887_406 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_407 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h197 == _T_481) begin
          _T_6887_407 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_408 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h198 == _T_481) begin
          _T_6887_408 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_409 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h199 == _T_481) begin
          _T_6887_409 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_410 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19a == _T_481) begin
          _T_6887_410 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_411 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19b == _T_481) begin
          _T_6887_411 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_412 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19c == _T_481) begin
          _T_6887_412 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_413 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19d == _T_481) begin
          _T_6887_413 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_414 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19e == _T_481) begin
          _T_6887_414 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_415 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h19f == _T_481) begin
          _T_6887_415 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_416 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a0 == _T_481) begin
          _T_6887_416 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_417 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a1 == _T_481) begin
          _T_6887_417 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_418 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a2 == _T_481) begin
          _T_6887_418 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_419 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a3 == _T_481) begin
          _T_6887_419 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_420 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a4 == _T_481) begin
          _T_6887_420 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_421 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a5 == _T_481) begin
          _T_6887_421 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_422 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a6 == _T_481) begin
          _T_6887_422 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_423 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a7 == _T_481) begin
          _T_6887_423 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_424 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a8 == _T_481) begin
          _T_6887_424 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_425 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1a9 == _T_481) begin
          _T_6887_425 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_426 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1aa == _T_481) begin
          _T_6887_426 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_427 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ab == _T_481) begin
          _T_6887_427 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_428 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ac == _T_481) begin
          _T_6887_428 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_429 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ad == _T_481) begin
          _T_6887_429 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_430 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ae == _T_481) begin
          _T_6887_430 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_431 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1af == _T_481) begin
          _T_6887_431 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_432 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b0 == _T_481) begin
          _T_6887_432 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_433 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b1 == _T_481) begin
          _T_6887_433 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_434 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b2 == _T_481) begin
          _T_6887_434 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_435 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b3 == _T_481) begin
          _T_6887_435 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_436 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b4 == _T_481) begin
          _T_6887_436 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_437 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b5 == _T_481) begin
          _T_6887_437 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_438 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b6 == _T_481) begin
          _T_6887_438 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_439 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b7 == _T_481) begin
          _T_6887_439 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_440 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b8 == _T_481) begin
          _T_6887_440 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_441 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1b9 == _T_481) begin
          _T_6887_441 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_442 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ba == _T_481) begin
          _T_6887_442 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_443 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1bb == _T_481) begin
          _T_6887_443 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_444 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1bc == _T_481) begin
          _T_6887_444 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_445 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1bd == _T_481) begin
          _T_6887_445 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_446 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1be == _T_481) begin
          _T_6887_446 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_447 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1bf == _T_481) begin
          _T_6887_447 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_448 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c0 == _T_481) begin
          _T_6887_448 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_449 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c1 == _T_481) begin
          _T_6887_449 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_450 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c2 == _T_481) begin
          _T_6887_450 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_451 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c3 == _T_481) begin
          _T_6887_451 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_452 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c4 == _T_481) begin
          _T_6887_452 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_453 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c5 == _T_481) begin
          _T_6887_453 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_454 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c6 == _T_481) begin
          _T_6887_454 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_455 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c7 == _T_481) begin
          _T_6887_455 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_456 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c8 == _T_481) begin
          _T_6887_456 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_457 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1c9 == _T_481) begin
          _T_6887_457 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_458 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ca == _T_481) begin
          _T_6887_458 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_459 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1cb == _T_481) begin
          _T_6887_459 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_460 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1cc == _T_481) begin
          _T_6887_460 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_461 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1cd == _T_481) begin
          _T_6887_461 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_462 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ce == _T_481) begin
          _T_6887_462 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_463 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1cf == _T_481) begin
          _T_6887_463 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_464 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d0 == _T_481) begin
          _T_6887_464 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_465 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d1 == _T_481) begin
          _T_6887_465 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_466 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d2 == _T_481) begin
          _T_6887_466 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_467 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d3 == _T_481) begin
          _T_6887_467 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_468 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d4 == _T_481) begin
          _T_6887_468 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_469 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d5 == _T_481) begin
          _T_6887_469 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_470 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d6 == _T_481) begin
          _T_6887_470 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_471 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d7 == _T_481) begin
          _T_6887_471 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_472 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d8 == _T_481) begin
          _T_6887_472 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_473 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1d9 == _T_481) begin
          _T_6887_473 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_474 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1da == _T_481) begin
          _T_6887_474 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_475 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1db == _T_481) begin
          _T_6887_475 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_476 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1dc == _T_481) begin
          _T_6887_476 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_477 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1dd == _T_481) begin
          _T_6887_477 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_478 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1de == _T_481) begin
          _T_6887_478 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_479 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1df == _T_481) begin
          _T_6887_479 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_480 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e0 == _T_481) begin
          _T_6887_480 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_481 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e1 == _T_481) begin
          _T_6887_481 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_482 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e2 == _T_481) begin
          _T_6887_482 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_483 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e3 == _T_481) begin
          _T_6887_483 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_484 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e4 == _T_481) begin
          _T_6887_484 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_485 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e5 == _T_481) begin
          _T_6887_485 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_486 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e6 == _T_481) begin
          _T_6887_486 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_487 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e7 == _T_481) begin
          _T_6887_487 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_488 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e8 == _T_481) begin
          _T_6887_488 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_489 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1e9 == _T_481) begin
          _T_6887_489 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_490 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ea == _T_481) begin
          _T_6887_490 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_491 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1eb == _T_481) begin
          _T_6887_491 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_492 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ec == _T_481) begin
          _T_6887_492 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_493 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ed == _T_481) begin
          _T_6887_493 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_494 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ee == _T_481) begin
          _T_6887_494 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_495 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ef == _T_481) begin
          _T_6887_495 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_496 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f0 == _T_481) begin
          _T_6887_496 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_497 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f1 == _T_481) begin
          _T_6887_497 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_498 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f2 == _T_481) begin
          _T_6887_498 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_499 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f3 == _T_481) begin
          _T_6887_499 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_500 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f4 == _T_481) begin
          _T_6887_500 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_501 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f5 == _T_481) begin
          _T_6887_501 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_502 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f6 == _T_481) begin
          _T_6887_502 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_503 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f7 == _T_481) begin
          _T_6887_503 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_504 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f8 == _T_481) begin
          _T_6887_504 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_505 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1f9 == _T_481) begin
          _T_6887_505 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_506 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1fa == _T_481) begin
          _T_6887_506 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_507 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1fb == _T_481) begin
          _T_6887_507 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_508 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1fc == _T_481) begin
          _T_6887_508 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_509 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1fd == _T_481) begin
          _T_6887_509 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_510 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1fe == _T_481) begin
          _T_6887_510 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_511 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h1ff == _T_481) begin
          _T_6887_511 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_512 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h200 == _T_481) begin
          _T_6887_512 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_513 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h201 == _T_481) begin
          _T_6887_513 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_514 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h202 == _T_481) begin
          _T_6887_514 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_515 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h203 == _T_481) begin
          _T_6887_515 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_516 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h204 == _T_481) begin
          _T_6887_516 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_517 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h205 == _T_481) begin
          _T_6887_517 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_518 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h206 == _T_481) begin
          _T_6887_518 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_519 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h207 == _T_481) begin
          _T_6887_519 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_520 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h208 == _T_481) begin
          _T_6887_520 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_521 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h209 == _T_481) begin
          _T_6887_521 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_522 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20a == _T_481) begin
          _T_6887_522 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_523 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20b == _T_481) begin
          _T_6887_523 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_524 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20c == _T_481) begin
          _T_6887_524 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_525 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20d == _T_481) begin
          _T_6887_525 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_526 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20e == _T_481) begin
          _T_6887_526 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_527 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h20f == _T_481) begin
          _T_6887_527 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_528 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h210 == _T_481) begin
          _T_6887_528 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_529 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h211 == _T_481) begin
          _T_6887_529 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_530 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h212 == _T_481) begin
          _T_6887_530 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_531 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h213 == _T_481) begin
          _T_6887_531 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_532 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h214 == _T_481) begin
          _T_6887_532 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_533 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h215 == _T_481) begin
          _T_6887_533 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_534 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h216 == _T_481) begin
          _T_6887_534 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_535 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h217 == _T_481) begin
          _T_6887_535 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_536 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h218 == _T_481) begin
          _T_6887_536 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_537 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h219 == _T_481) begin
          _T_6887_537 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_538 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21a == _T_481) begin
          _T_6887_538 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_539 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21b == _T_481) begin
          _T_6887_539 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_540 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21c == _T_481) begin
          _T_6887_540 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_541 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21d == _T_481) begin
          _T_6887_541 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_542 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21e == _T_481) begin
          _T_6887_542 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_543 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h21f == _T_481) begin
          _T_6887_543 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_544 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h220 == _T_481) begin
          _T_6887_544 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_545 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h221 == _T_481) begin
          _T_6887_545 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_546 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h222 == _T_481) begin
          _T_6887_546 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_547 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h223 == _T_481) begin
          _T_6887_547 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_548 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h224 == _T_481) begin
          _T_6887_548 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_549 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h225 == _T_481) begin
          _T_6887_549 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_550 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h226 == _T_481) begin
          _T_6887_550 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_551 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h227 == _T_481) begin
          _T_6887_551 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_552 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h228 == _T_481) begin
          _T_6887_552 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_553 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h229 == _T_481) begin
          _T_6887_553 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_554 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22a == _T_481) begin
          _T_6887_554 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_555 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22b == _T_481) begin
          _T_6887_555 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_556 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22c == _T_481) begin
          _T_6887_556 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_557 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22d == _T_481) begin
          _T_6887_557 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_558 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22e == _T_481) begin
          _T_6887_558 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_559 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h22f == _T_481) begin
          _T_6887_559 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_560 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h230 == _T_481) begin
          _T_6887_560 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_561 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h231 == _T_481) begin
          _T_6887_561 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_562 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h232 == _T_481) begin
          _T_6887_562 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_563 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h233 == _T_481) begin
          _T_6887_563 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_564 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h234 == _T_481) begin
          _T_6887_564 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_565 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h235 == _T_481) begin
          _T_6887_565 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_566 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h236 == _T_481) begin
          _T_6887_566 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_567 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h237 == _T_481) begin
          _T_6887_567 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_568 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h238 == _T_481) begin
          _T_6887_568 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_569 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h239 == _T_481) begin
          _T_6887_569 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_570 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23a == _T_481) begin
          _T_6887_570 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_571 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23b == _T_481) begin
          _T_6887_571 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_572 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23c == _T_481) begin
          _T_6887_572 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_573 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23d == _T_481) begin
          _T_6887_573 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_574 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23e == _T_481) begin
          _T_6887_574 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_575 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h23f == _T_481) begin
          _T_6887_575 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_576 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h240 == _T_481) begin
          _T_6887_576 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_577 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h241 == _T_481) begin
          _T_6887_577 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_578 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h242 == _T_481) begin
          _T_6887_578 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_579 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h243 == _T_481) begin
          _T_6887_579 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_580 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h244 == _T_481) begin
          _T_6887_580 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_581 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h245 == _T_481) begin
          _T_6887_581 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_582 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h246 == _T_481) begin
          _T_6887_582 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_583 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h247 == _T_481) begin
          _T_6887_583 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_584 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h248 == _T_481) begin
          _T_6887_584 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_585 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h249 == _T_481) begin
          _T_6887_585 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_586 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24a == _T_481) begin
          _T_6887_586 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_587 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24b == _T_481) begin
          _T_6887_587 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_588 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24c == _T_481) begin
          _T_6887_588 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_589 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24d == _T_481) begin
          _T_6887_589 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_590 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24e == _T_481) begin
          _T_6887_590 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_591 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h24f == _T_481) begin
          _T_6887_591 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_592 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h250 == _T_481) begin
          _T_6887_592 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_593 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h251 == _T_481) begin
          _T_6887_593 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_594 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h252 == _T_481) begin
          _T_6887_594 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_595 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h253 == _T_481) begin
          _T_6887_595 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_596 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h254 == _T_481) begin
          _T_6887_596 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_597 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h255 == _T_481) begin
          _T_6887_597 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_598 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h256 == _T_481) begin
          _T_6887_598 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_599 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h257 == _T_481) begin
          _T_6887_599 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_600 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h258 == _T_481) begin
          _T_6887_600 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_601 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h259 == _T_481) begin
          _T_6887_601 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_602 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25a == _T_481) begin
          _T_6887_602 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_603 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25b == _T_481) begin
          _T_6887_603 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_604 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25c == _T_481) begin
          _T_6887_604 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_605 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25d == _T_481) begin
          _T_6887_605 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_606 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25e == _T_481) begin
          _T_6887_606 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_607 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h25f == _T_481) begin
          _T_6887_607 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_608 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h260 == _T_481) begin
          _T_6887_608 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_609 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h261 == _T_481) begin
          _T_6887_609 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_610 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h262 == _T_481) begin
          _T_6887_610 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_611 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h263 == _T_481) begin
          _T_6887_611 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_612 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h264 == _T_481) begin
          _T_6887_612 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_613 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h265 == _T_481) begin
          _T_6887_613 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_614 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h266 == _T_481) begin
          _T_6887_614 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_615 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h267 == _T_481) begin
          _T_6887_615 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_616 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h268 == _T_481) begin
          _T_6887_616 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_617 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h269 == _T_481) begin
          _T_6887_617 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_618 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26a == _T_481) begin
          _T_6887_618 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_619 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26b == _T_481) begin
          _T_6887_619 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_620 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26c == _T_481) begin
          _T_6887_620 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_621 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26d == _T_481) begin
          _T_6887_621 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_622 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26e == _T_481) begin
          _T_6887_622 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_623 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h26f == _T_481) begin
          _T_6887_623 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_624 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h270 == _T_481) begin
          _T_6887_624 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_625 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h271 == _T_481) begin
          _T_6887_625 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_626 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h272 == _T_481) begin
          _T_6887_626 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_627 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h273 == _T_481) begin
          _T_6887_627 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_628 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h274 == _T_481) begin
          _T_6887_628 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_629 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h275 == _T_481) begin
          _T_6887_629 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_630 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h276 == _T_481) begin
          _T_6887_630 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_631 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h277 == _T_481) begin
          _T_6887_631 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_632 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h278 == _T_481) begin
          _T_6887_632 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_633 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h279 == _T_481) begin
          _T_6887_633 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_634 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27a == _T_481) begin
          _T_6887_634 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_635 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27b == _T_481) begin
          _T_6887_635 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_636 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27c == _T_481) begin
          _T_6887_636 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_637 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27d == _T_481) begin
          _T_6887_637 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_638 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27e == _T_481) begin
          _T_6887_638 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_639 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h27f == _T_481) begin
          _T_6887_639 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_640 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h280 == _T_481) begin
          _T_6887_640 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_641 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h281 == _T_481) begin
          _T_6887_641 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_642 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h282 == _T_481) begin
          _T_6887_642 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_643 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h283 == _T_481) begin
          _T_6887_643 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_644 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h284 == _T_481) begin
          _T_6887_644 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_645 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h285 == _T_481) begin
          _T_6887_645 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_646 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h286 == _T_481) begin
          _T_6887_646 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_647 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h287 == _T_481) begin
          _T_6887_647 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_648 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h288 == _T_481) begin
          _T_6887_648 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_649 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h289 == _T_481) begin
          _T_6887_649 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_650 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28a == _T_481) begin
          _T_6887_650 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_651 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28b == _T_481) begin
          _T_6887_651 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_652 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28c == _T_481) begin
          _T_6887_652 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_653 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28d == _T_481) begin
          _T_6887_653 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_654 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28e == _T_481) begin
          _T_6887_654 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_655 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h28f == _T_481) begin
          _T_6887_655 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_656 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h290 == _T_481) begin
          _T_6887_656 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_657 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h291 == _T_481) begin
          _T_6887_657 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_658 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h292 == _T_481) begin
          _T_6887_658 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_659 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h293 == _T_481) begin
          _T_6887_659 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_660 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h294 == _T_481) begin
          _T_6887_660 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_661 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h295 == _T_481) begin
          _T_6887_661 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_662 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h296 == _T_481) begin
          _T_6887_662 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_663 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h297 == _T_481) begin
          _T_6887_663 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_664 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h298 == _T_481) begin
          _T_6887_664 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_665 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h299 == _T_481) begin
          _T_6887_665 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_666 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29a == _T_481) begin
          _T_6887_666 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_667 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29b == _T_481) begin
          _T_6887_667 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_668 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29c == _T_481) begin
          _T_6887_668 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_669 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29d == _T_481) begin
          _T_6887_669 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_670 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29e == _T_481) begin
          _T_6887_670 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_671 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h29f == _T_481) begin
          _T_6887_671 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_672 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a0 == _T_481) begin
          _T_6887_672 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_673 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a1 == _T_481) begin
          _T_6887_673 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_674 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a2 == _T_481) begin
          _T_6887_674 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_675 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a3 == _T_481) begin
          _T_6887_675 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_676 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a4 == _T_481) begin
          _T_6887_676 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_677 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a5 == _T_481) begin
          _T_6887_677 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_678 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a6 == _T_481) begin
          _T_6887_678 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_679 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a7 == _T_481) begin
          _T_6887_679 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_680 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a8 == _T_481) begin
          _T_6887_680 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_681 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2a9 == _T_481) begin
          _T_6887_681 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_682 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2aa == _T_481) begin
          _T_6887_682 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_683 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ab == _T_481) begin
          _T_6887_683 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_684 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ac == _T_481) begin
          _T_6887_684 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_685 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ad == _T_481) begin
          _T_6887_685 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_686 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ae == _T_481) begin
          _T_6887_686 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_687 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2af == _T_481) begin
          _T_6887_687 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_688 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b0 == _T_481) begin
          _T_6887_688 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_689 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b1 == _T_481) begin
          _T_6887_689 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_690 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b2 == _T_481) begin
          _T_6887_690 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_691 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b3 == _T_481) begin
          _T_6887_691 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_692 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b4 == _T_481) begin
          _T_6887_692 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_693 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b5 == _T_481) begin
          _T_6887_693 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_694 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b6 == _T_481) begin
          _T_6887_694 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_695 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b7 == _T_481) begin
          _T_6887_695 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_696 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b8 == _T_481) begin
          _T_6887_696 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_697 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2b9 == _T_481) begin
          _T_6887_697 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_698 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ba == _T_481) begin
          _T_6887_698 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_699 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2bb == _T_481) begin
          _T_6887_699 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_700 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2bc == _T_481) begin
          _T_6887_700 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_701 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2bd == _T_481) begin
          _T_6887_701 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_702 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2be == _T_481) begin
          _T_6887_702 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_703 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2bf == _T_481) begin
          _T_6887_703 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_704 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c0 == _T_481) begin
          _T_6887_704 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_705 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c1 == _T_481) begin
          _T_6887_705 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_706 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c2 == _T_481) begin
          _T_6887_706 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_707 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c3 == _T_481) begin
          _T_6887_707 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_708 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c4 == _T_481) begin
          _T_6887_708 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_709 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c5 == _T_481) begin
          _T_6887_709 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_710 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c6 == _T_481) begin
          _T_6887_710 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_711 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c7 == _T_481) begin
          _T_6887_711 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_712 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c8 == _T_481) begin
          _T_6887_712 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_713 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2c9 == _T_481) begin
          _T_6887_713 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_714 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ca == _T_481) begin
          _T_6887_714 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_715 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2cb == _T_481) begin
          _T_6887_715 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_716 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2cc == _T_481) begin
          _T_6887_716 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_717 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2cd == _T_481) begin
          _T_6887_717 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_718 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ce == _T_481) begin
          _T_6887_718 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_719 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2cf == _T_481) begin
          _T_6887_719 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_720 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d0 == _T_481) begin
          _T_6887_720 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_721 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d1 == _T_481) begin
          _T_6887_721 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_722 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d2 == _T_481) begin
          _T_6887_722 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_723 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d3 == _T_481) begin
          _T_6887_723 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_724 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d4 == _T_481) begin
          _T_6887_724 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_725 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d5 == _T_481) begin
          _T_6887_725 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_726 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d6 == _T_481) begin
          _T_6887_726 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_727 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d7 == _T_481) begin
          _T_6887_727 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_728 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d8 == _T_481) begin
          _T_6887_728 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_729 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2d9 == _T_481) begin
          _T_6887_729 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_730 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2da == _T_481) begin
          _T_6887_730 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_731 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2db == _T_481) begin
          _T_6887_731 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_732 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2dc == _T_481) begin
          _T_6887_732 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_733 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2dd == _T_481) begin
          _T_6887_733 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_734 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2de == _T_481) begin
          _T_6887_734 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_735 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2df == _T_481) begin
          _T_6887_735 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_736 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e0 == _T_481) begin
          _T_6887_736 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_737 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e1 == _T_481) begin
          _T_6887_737 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_738 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e2 == _T_481) begin
          _T_6887_738 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_739 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e3 == _T_481) begin
          _T_6887_739 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_740 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e4 == _T_481) begin
          _T_6887_740 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_741 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e5 == _T_481) begin
          _T_6887_741 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_742 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e6 == _T_481) begin
          _T_6887_742 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_743 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e7 == _T_481) begin
          _T_6887_743 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_744 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e8 == _T_481) begin
          _T_6887_744 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_745 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2e9 == _T_481) begin
          _T_6887_745 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_746 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ea == _T_481) begin
          _T_6887_746 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_747 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2eb == _T_481) begin
          _T_6887_747 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_748 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ec == _T_481) begin
          _T_6887_748 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_749 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ed == _T_481) begin
          _T_6887_749 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_750 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ee == _T_481) begin
          _T_6887_750 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_751 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ef == _T_481) begin
          _T_6887_751 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_752 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f0 == _T_481) begin
          _T_6887_752 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_753 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f1 == _T_481) begin
          _T_6887_753 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_754 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f2 == _T_481) begin
          _T_6887_754 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_755 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f3 == _T_481) begin
          _T_6887_755 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_756 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f4 == _T_481) begin
          _T_6887_756 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_757 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f5 == _T_481) begin
          _T_6887_757 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_758 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f6 == _T_481) begin
          _T_6887_758 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_759 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f7 == _T_481) begin
          _T_6887_759 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_760 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f8 == _T_481) begin
          _T_6887_760 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_761 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2f9 == _T_481) begin
          _T_6887_761 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_762 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2fa == _T_481) begin
          _T_6887_762 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_763 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2fb == _T_481) begin
          _T_6887_763 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_764 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2fc == _T_481) begin
          _T_6887_764 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_765 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2fd == _T_481) begin
          _T_6887_765 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_766 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2fe == _T_481) begin
          _T_6887_766 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_767 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h2ff == _T_481) begin
          _T_6887_767 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_768 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h300 == _T_481) begin
          _T_6887_768 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_769 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h301 == _T_481) begin
          _T_6887_769 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_770 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h302 == _T_481) begin
          _T_6887_770 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_771 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h303 == _T_481) begin
          _T_6887_771 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_772 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h304 == _T_481) begin
          _T_6887_772 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_773 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h305 == _T_481) begin
          _T_6887_773 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_774 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h306 == _T_481) begin
          _T_6887_774 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_775 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h307 == _T_481) begin
          _T_6887_775 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_776 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h308 == _T_481) begin
          _T_6887_776 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_777 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h309 == _T_481) begin
          _T_6887_777 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_778 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30a == _T_481) begin
          _T_6887_778 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_779 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30b == _T_481) begin
          _T_6887_779 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_780 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30c == _T_481) begin
          _T_6887_780 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_781 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30d == _T_481) begin
          _T_6887_781 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_782 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30e == _T_481) begin
          _T_6887_782 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_783 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h30f == _T_481) begin
          _T_6887_783 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_784 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h310 == _T_481) begin
          _T_6887_784 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_785 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h311 == _T_481) begin
          _T_6887_785 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_786 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h312 == _T_481) begin
          _T_6887_786 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_787 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h313 == _T_481) begin
          _T_6887_787 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_788 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h314 == _T_481) begin
          _T_6887_788 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_789 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h315 == _T_481) begin
          _T_6887_789 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_790 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h316 == _T_481) begin
          _T_6887_790 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_791 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h317 == _T_481) begin
          _T_6887_791 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_792 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h318 == _T_481) begin
          _T_6887_792 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_793 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h319 == _T_481) begin
          _T_6887_793 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_794 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31a == _T_481) begin
          _T_6887_794 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_795 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31b == _T_481) begin
          _T_6887_795 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_796 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31c == _T_481) begin
          _T_6887_796 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_797 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31d == _T_481) begin
          _T_6887_797 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_798 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31e == _T_481) begin
          _T_6887_798 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_799 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h31f == _T_481) begin
          _T_6887_799 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_800 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h320 == _T_481) begin
          _T_6887_800 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_801 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h321 == _T_481) begin
          _T_6887_801 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_802 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h322 == _T_481) begin
          _T_6887_802 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_803 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h323 == _T_481) begin
          _T_6887_803 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_804 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h324 == _T_481) begin
          _T_6887_804 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_805 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h325 == _T_481) begin
          _T_6887_805 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_806 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h326 == _T_481) begin
          _T_6887_806 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_807 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h327 == _T_481) begin
          _T_6887_807 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_808 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h328 == _T_481) begin
          _T_6887_808 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_809 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h329 == _T_481) begin
          _T_6887_809 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_810 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32a == _T_481) begin
          _T_6887_810 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_811 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32b == _T_481) begin
          _T_6887_811 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_812 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32c == _T_481) begin
          _T_6887_812 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_813 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32d == _T_481) begin
          _T_6887_813 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_814 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32e == _T_481) begin
          _T_6887_814 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_815 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h32f == _T_481) begin
          _T_6887_815 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_816 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h330 == _T_481) begin
          _T_6887_816 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_817 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h331 == _T_481) begin
          _T_6887_817 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_818 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h332 == _T_481) begin
          _T_6887_818 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_819 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h333 == _T_481) begin
          _T_6887_819 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_820 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h334 == _T_481) begin
          _T_6887_820 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_821 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h335 == _T_481) begin
          _T_6887_821 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_822 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h336 == _T_481) begin
          _T_6887_822 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_823 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h337 == _T_481) begin
          _T_6887_823 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_824 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h338 == _T_481) begin
          _T_6887_824 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_825 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h339 == _T_481) begin
          _T_6887_825 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_826 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33a == _T_481) begin
          _T_6887_826 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_827 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33b == _T_481) begin
          _T_6887_827 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_828 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33c == _T_481) begin
          _T_6887_828 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_829 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33d == _T_481) begin
          _T_6887_829 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_830 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33e == _T_481) begin
          _T_6887_830 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_831 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h33f == _T_481) begin
          _T_6887_831 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_832 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h340 == _T_481) begin
          _T_6887_832 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_833 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h341 == _T_481) begin
          _T_6887_833 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_834 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h342 == _T_481) begin
          _T_6887_834 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_835 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h343 == _T_481) begin
          _T_6887_835 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_836 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h344 == _T_481) begin
          _T_6887_836 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_837 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h345 == _T_481) begin
          _T_6887_837 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_838 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h346 == _T_481) begin
          _T_6887_838 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_839 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h347 == _T_481) begin
          _T_6887_839 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_840 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h348 == _T_481) begin
          _T_6887_840 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_841 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h349 == _T_481) begin
          _T_6887_841 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_842 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34a == _T_481) begin
          _T_6887_842 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_843 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34b == _T_481) begin
          _T_6887_843 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_844 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34c == _T_481) begin
          _T_6887_844 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_845 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34d == _T_481) begin
          _T_6887_845 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_846 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34e == _T_481) begin
          _T_6887_846 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_847 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h34f == _T_481) begin
          _T_6887_847 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_848 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h350 == _T_481) begin
          _T_6887_848 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_849 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h351 == _T_481) begin
          _T_6887_849 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_850 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h352 == _T_481) begin
          _T_6887_850 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_851 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h353 == _T_481) begin
          _T_6887_851 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_852 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h354 == _T_481) begin
          _T_6887_852 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_853 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h355 == _T_481) begin
          _T_6887_853 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_854 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h356 == _T_481) begin
          _T_6887_854 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_855 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h357 == _T_481) begin
          _T_6887_855 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_856 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h358 == _T_481) begin
          _T_6887_856 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_857 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h359 == _T_481) begin
          _T_6887_857 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_858 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35a == _T_481) begin
          _T_6887_858 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_859 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35b == _T_481) begin
          _T_6887_859 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_860 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35c == _T_481) begin
          _T_6887_860 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_861 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35d == _T_481) begin
          _T_6887_861 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_862 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35e == _T_481) begin
          _T_6887_862 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_863 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h35f == _T_481) begin
          _T_6887_863 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_864 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h360 == _T_481) begin
          _T_6887_864 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_865 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h361 == _T_481) begin
          _T_6887_865 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_866 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h362 == _T_481) begin
          _T_6887_866 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_867 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h363 == _T_481) begin
          _T_6887_867 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_868 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h364 == _T_481) begin
          _T_6887_868 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_869 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h365 == _T_481) begin
          _T_6887_869 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_870 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h366 == _T_481) begin
          _T_6887_870 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_871 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h367 == _T_481) begin
          _T_6887_871 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_872 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h368 == _T_481) begin
          _T_6887_872 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_873 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h369 == _T_481) begin
          _T_6887_873 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_874 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36a == _T_481) begin
          _T_6887_874 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_875 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36b == _T_481) begin
          _T_6887_875 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_876 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36c == _T_481) begin
          _T_6887_876 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_877 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36d == _T_481) begin
          _T_6887_877 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_878 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36e == _T_481) begin
          _T_6887_878 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_879 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h36f == _T_481) begin
          _T_6887_879 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_880 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h370 == _T_481) begin
          _T_6887_880 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_881 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h371 == _T_481) begin
          _T_6887_881 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_882 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h372 == _T_481) begin
          _T_6887_882 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_883 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h373 == _T_481) begin
          _T_6887_883 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_884 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h374 == _T_481) begin
          _T_6887_884 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_885 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h375 == _T_481) begin
          _T_6887_885 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_886 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h376 == _T_481) begin
          _T_6887_886 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_887 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h377 == _T_481) begin
          _T_6887_887 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_888 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h378 == _T_481) begin
          _T_6887_888 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_889 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h379 == _T_481) begin
          _T_6887_889 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_890 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37a == _T_481) begin
          _T_6887_890 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_891 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37b == _T_481) begin
          _T_6887_891 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_892 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37c == _T_481) begin
          _T_6887_892 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_893 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37d == _T_481) begin
          _T_6887_893 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_894 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37e == _T_481) begin
          _T_6887_894 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_895 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h37f == _T_481) begin
          _T_6887_895 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_896 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h380 == _T_481) begin
          _T_6887_896 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_897 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h381 == _T_481) begin
          _T_6887_897 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_898 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h382 == _T_481) begin
          _T_6887_898 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_899 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h383 == _T_481) begin
          _T_6887_899 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_900 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h384 == _T_481) begin
          _T_6887_900 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_901 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h385 == _T_481) begin
          _T_6887_901 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_902 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h386 == _T_481) begin
          _T_6887_902 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_903 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h387 == _T_481) begin
          _T_6887_903 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_904 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h388 == _T_481) begin
          _T_6887_904 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_905 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h389 == _T_481) begin
          _T_6887_905 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_906 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38a == _T_481) begin
          _T_6887_906 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_907 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38b == _T_481) begin
          _T_6887_907 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_908 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38c == _T_481) begin
          _T_6887_908 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_909 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38d == _T_481) begin
          _T_6887_909 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_910 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38e == _T_481) begin
          _T_6887_910 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_911 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h38f == _T_481) begin
          _T_6887_911 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_912 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h390 == _T_481) begin
          _T_6887_912 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_913 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h391 == _T_481) begin
          _T_6887_913 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_914 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h392 == _T_481) begin
          _T_6887_914 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_915 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h393 == _T_481) begin
          _T_6887_915 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_916 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h394 == _T_481) begin
          _T_6887_916 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_917 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h395 == _T_481) begin
          _T_6887_917 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_918 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h396 == _T_481) begin
          _T_6887_918 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_919 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h397 == _T_481) begin
          _T_6887_919 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_920 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h398 == _T_481) begin
          _T_6887_920 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_921 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h399 == _T_481) begin
          _T_6887_921 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_922 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39a == _T_481) begin
          _T_6887_922 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_923 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39b == _T_481) begin
          _T_6887_923 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_924 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39c == _T_481) begin
          _T_6887_924 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_925 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39d == _T_481) begin
          _T_6887_925 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_926 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39e == _T_481) begin
          _T_6887_926 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_927 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h39f == _T_481) begin
          _T_6887_927 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_928 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a0 == _T_481) begin
          _T_6887_928 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_929 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a1 == _T_481) begin
          _T_6887_929 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_930 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a2 == _T_481) begin
          _T_6887_930 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_931 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a3 == _T_481) begin
          _T_6887_931 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_932 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a4 == _T_481) begin
          _T_6887_932 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_933 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a5 == _T_481) begin
          _T_6887_933 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_934 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a6 == _T_481) begin
          _T_6887_934 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_935 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a7 == _T_481) begin
          _T_6887_935 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_936 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a8 == _T_481) begin
          _T_6887_936 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_937 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3a9 == _T_481) begin
          _T_6887_937 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_938 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3aa == _T_481) begin
          _T_6887_938 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_939 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ab == _T_481) begin
          _T_6887_939 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_940 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ac == _T_481) begin
          _T_6887_940 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_941 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ad == _T_481) begin
          _T_6887_941 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_942 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ae == _T_481) begin
          _T_6887_942 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_943 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3af == _T_481) begin
          _T_6887_943 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_944 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b0 == _T_481) begin
          _T_6887_944 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_945 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b1 == _T_481) begin
          _T_6887_945 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_946 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b2 == _T_481) begin
          _T_6887_946 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_947 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b3 == _T_481) begin
          _T_6887_947 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_948 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b4 == _T_481) begin
          _T_6887_948 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_949 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b5 == _T_481) begin
          _T_6887_949 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_950 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b6 == _T_481) begin
          _T_6887_950 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_951 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b7 == _T_481) begin
          _T_6887_951 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_952 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b8 == _T_481) begin
          _T_6887_952 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_953 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3b9 == _T_481) begin
          _T_6887_953 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_954 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ba == _T_481) begin
          _T_6887_954 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_955 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3bb == _T_481) begin
          _T_6887_955 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_956 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3bc == _T_481) begin
          _T_6887_956 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_957 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3bd == _T_481) begin
          _T_6887_957 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_958 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3be == _T_481) begin
          _T_6887_958 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_959 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3bf == _T_481) begin
          _T_6887_959 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_960 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c0 == _T_481) begin
          _T_6887_960 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_961 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c1 == _T_481) begin
          _T_6887_961 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_962 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c2 == _T_481) begin
          _T_6887_962 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_963 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c3 == _T_481) begin
          _T_6887_963 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_964 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c4 == _T_481) begin
          _T_6887_964 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_965 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c5 == _T_481) begin
          _T_6887_965 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_966 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c6 == _T_481) begin
          _T_6887_966 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_967 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c7 == _T_481) begin
          _T_6887_967 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_968 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c8 == _T_481) begin
          _T_6887_968 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_969 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3c9 == _T_481) begin
          _T_6887_969 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_970 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ca == _T_481) begin
          _T_6887_970 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_971 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3cb == _T_481) begin
          _T_6887_971 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_972 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3cc == _T_481) begin
          _T_6887_972 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_973 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3cd == _T_481) begin
          _T_6887_973 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_974 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ce == _T_481) begin
          _T_6887_974 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_975 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3cf == _T_481) begin
          _T_6887_975 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_976 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d0 == _T_481) begin
          _T_6887_976 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_977 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d1 == _T_481) begin
          _T_6887_977 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_978 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d2 == _T_481) begin
          _T_6887_978 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_979 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d3 == _T_481) begin
          _T_6887_979 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_980 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d4 == _T_481) begin
          _T_6887_980 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_981 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d5 == _T_481) begin
          _T_6887_981 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_982 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d6 == _T_481) begin
          _T_6887_982 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_983 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d7 == _T_481) begin
          _T_6887_983 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_984 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d8 == _T_481) begin
          _T_6887_984 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_985 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3d9 == _T_481) begin
          _T_6887_985 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_986 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3da == _T_481) begin
          _T_6887_986 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_987 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3db == _T_481) begin
          _T_6887_987 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_988 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3dc == _T_481) begin
          _T_6887_988 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_989 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3dd == _T_481) begin
          _T_6887_989 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_990 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3de == _T_481) begin
          _T_6887_990 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_991 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3df == _T_481) begin
          _T_6887_991 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_992 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e0 == _T_481) begin
          _T_6887_992 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_993 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e1 == _T_481) begin
          _T_6887_993 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_994 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e2 == _T_481) begin
          _T_6887_994 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_995 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e3 == _T_481) begin
          _T_6887_995 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_996 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e4 == _T_481) begin
          _T_6887_996 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_997 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e5 == _T_481) begin
          _T_6887_997 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_998 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e6 == _T_481) begin
          _T_6887_998 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_999 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e7 == _T_481) begin
          _T_6887_999 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1000 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e8 == _T_481) begin
          _T_6887_1000 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1001 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3e9 == _T_481) begin
          _T_6887_1001 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1002 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ea == _T_481) begin
          _T_6887_1002 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1003 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3eb == _T_481) begin
          _T_6887_1003 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1004 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ec == _T_481) begin
          _T_6887_1004 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1005 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ed == _T_481) begin
          _T_6887_1005 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1006 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ee == _T_481) begin
          _T_6887_1006 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1007 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ef == _T_481) begin
          _T_6887_1007 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1008 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f0 == _T_481) begin
          _T_6887_1008 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1009 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f1 == _T_481) begin
          _T_6887_1009 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1010 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f2 == _T_481) begin
          _T_6887_1010 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1011 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f3 == _T_481) begin
          _T_6887_1011 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1012 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f4 == _T_481) begin
          _T_6887_1012 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1013 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f5 == _T_481) begin
          _T_6887_1013 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1014 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f6 == _T_481) begin
          _T_6887_1014 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1015 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f7 == _T_481) begin
          _T_6887_1015 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1016 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f8 == _T_481) begin
          _T_6887_1016 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1017 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3f9 == _T_481) begin
          _T_6887_1017 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1018 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3fa == _T_481) begin
          _T_6887_1018 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1019 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3fb == _T_481) begin
          _T_6887_1019 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1020 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3fc == _T_481) begin
          _T_6887_1020 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1021 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3fd == _T_481) begin
          _T_6887_1021 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1022 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3fe == _T_481) begin
          _T_6887_1022 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1023 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h3ff == _T_481) begin
          _T_6887_1023 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1024 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h400 == _T_481) begin
          _T_6887_1024 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1025 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h401 == _T_481) begin
          _T_6887_1025 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1026 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h402 == _T_481) begin
          _T_6887_1026 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1027 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h403 == _T_481) begin
          _T_6887_1027 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1028 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h404 == _T_481) begin
          _T_6887_1028 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1029 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h405 == _T_481) begin
          _T_6887_1029 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1030 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h406 == _T_481) begin
          _T_6887_1030 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1031 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h407 == _T_481) begin
          _T_6887_1031 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1032 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h408 == _T_481) begin
          _T_6887_1032 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1033 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h409 == _T_481) begin
          _T_6887_1033 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1034 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40a == _T_481) begin
          _T_6887_1034 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1035 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40b == _T_481) begin
          _T_6887_1035 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1036 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40c == _T_481) begin
          _T_6887_1036 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1037 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40d == _T_481) begin
          _T_6887_1037 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1038 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40e == _T_481) begin
          _T_6887_1038 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1039 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h40f == _T_481) begin
          _T_6887_1039 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1040 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h410 == _T_481) begin
          _T_6887_1040 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1041 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h411 == _T_481) begin
          _T_6887_1041 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1042 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h412 == _T_481) begin
          _T_6887_1042 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1043 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h413 == _T_481) begin
          _T_6887_1043 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1044 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h414 == _T_481) begin
          _T_6887_1044 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1045 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h415 == _T_481) begin
          _T_6887_1045 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1046 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h416 == _T_481) begin
          _T_6887_1046 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1047 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h417 == _T_481) begin
          _T_6887_1047 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1048 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h418 == _T_481) begin
          _T_6887_1048 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1049 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h419 == _T_481) begin
          _T_6887_1049 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1050 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41a == _T_481) begin
          _T_6887_1050 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1051 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41b == _T_481) begin
          _T_6887_1051 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1052 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41c == _T_481) begin
          _T_6887_1052 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1053 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41d == _T_481) begin
          _T_6887_1053 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1054 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41e == _T_481) begin
          _T_6887_1054 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1055 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h41f == _T_481) begin
          _T_6887_1055 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1056 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h420 == _T_481) begin
          _T_6887_1056 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1057 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h421 == _T_481) begin
          _T_6887_1057 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1058 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h422 == _T_481) begin
          _T_6887_1058 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1059 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h423 == _T_481) begin
          _T_6887_1059 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1060 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h424 == _T_481) begin
          _T_6887_1060 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1061 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h425 == _T_481) begin
          _T_6887_1061 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1062 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h426 == _T_481) begin
          _T_6887_1062 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1063 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h427 == _T_481) begin
          _T_6887_1063 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1064 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h428 == _T_481) begin
          _T_6887_1064 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1065 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h429 == _T_481) begin
          _T_6887_1065 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1066 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42a == _T_481) begin
          _T_6887_1066 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1067 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42b == _T_481) begin
          _T_6887_1067 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1068 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42c == _T_481) begin
          _T_6887_1068 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1069 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42d == _T_481) begin
          _T_6887_1069 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1070 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42e == _T_481) begin
          _T_6887_1070 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1071 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h42f == _T_481) begin
          _T_6887_1071 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1072 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h430 == _T_481) begin
          _T_6887_1072 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1073 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h431 == _T_481) begin
          _T_6887_1073 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1074 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h432 == _T_481) begin
          _T_6887_1074 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1075 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h433 == _T_481) begin
          _T_6887_1075 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1076 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h434 == _T_481) begin
          _T_6887_1076 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1077 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h435 == _T_481) begin
          _T_6887_1077 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1078 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h436 == _T_481) begin
          _T_6887_1078 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1079 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h437 == _T_481) begin
          _T_6887_1079 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1080 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h438 == _T_481) begin
          _T_6887_1080 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1081 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h439 == _T_481) begin
          _T_6887_1081 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1082 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43a == _T_481) begin
          _T_6887_1082 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1083 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43b == _T_481) begin
          _T_6887_1083 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1084 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43c == _T_481) begin
          _T_6887_1084 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1085 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43d == _T_481) begin
          _T_6887_1085 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1086 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43e == _T_481) begin
          _T_6887_1086 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1087 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h43f == _T_481) begin
          _T_6887_1087 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1088 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h440 == _T_481) begin
          _T_6887_1088 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1089 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h441 == _T_481) begin
          _T_6887_1089 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1090 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h442 == _T_481) begin
          _T_6887_1090 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1091 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h443 == _T_481) begin
          _T_6887_1091 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1092 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h444 == _T_481) begin
          _T_6887_1092 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1093 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h445 == _T_481) begin
          _T_6887_1093 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1094 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h446 == _T_481) begin
          _T_6887_1094 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1095 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h447 == _T_481) begin
          _T_6887_1095 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1096 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h448 == _T_481) begin
          _T_6887_1096 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1097 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h449 == _T_481) begin
          _T_6887_1097 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1098 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44a == _T_481) begin
          _T_6887_1098 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1099 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44b == _T_481) begin
          _T_6887_1099 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1100 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44c == _T_481) begin
          _T_6887_1100 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1101 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44d == _T_481) begin
          _T_6887_1101 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1102 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44e == _T_481) begin
          _T_6887_1102 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1103 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h44f == _T_481) begin
          _T_6887_1103 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1104 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h450 == _T_481) begin
          _T_6887_1104 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1105 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h451 == _T_481) begin
          _T_6887_1105 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1106 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h452 == _T_481) begin
          _T_6887_1106 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1107 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h453 == _T_481) begin
          _T_6887_1107 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1108 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h454 == _T_481) begin
          _T_6887_1108 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1109 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h455 == _T_481) begin
          _T_6887_1109 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1110 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h456 == _T_481) begin
          _T_6887_1110 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1111 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h457 == _T_481) begin
          _T_6887_1111 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1112 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h458 == _T_481) begin
          _T_6887_1112 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1113 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h459 == _T_481) begin
          _T_6887_1113 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1114 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45a == _T_481) begin
          _T_6887_1114 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1115 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45b == _T_481) begin
          _T_6887_1115 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1116 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45c == _T_481) begin
          _T_6887_1116 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1117 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45d == _T_481) begin
          _T_6887_1117 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1118 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45e == _T_481) begin
          _T_6887_1118 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1119 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h45f == _T_481) begin
          _T_6887_1119 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1120 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h460 == _T_481) begin
          _T_6887_1120 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1121 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h461 == _T_481) begin
          _T_6887_1121 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1122 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h462 == _T_481) begin
          _T_6887_1122 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1123 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h463 == _T_481) begin
          _T_6887_1123 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1124 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h464 == _T_481) begin
          _T_6887_1124 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1125 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h465 == _T_481) begin
          _T_6887_1125 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1126 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h466 == _T_481) begin
          _T_6887_1126 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1127 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h467 == _T_481) begin
          _T_6887_1127 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1128 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h468 == _T_481) begin
          _T_6887_1128 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1129 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h469 == _T_481) begin
          _T_6887_1129 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1130 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46a == _T_481) begin
          _T_6887_1130 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1131 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46b == _T_481) begin
          _T_6887_1131 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1132 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46c == _T_481) begin
          _T_6887_1132 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1133 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46d == _T_481) begin
          _T_6887_1133 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1134 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46e == _T_481) begin
          _T_6887_1134 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1135 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h46f == _T_481) begin
          _T_6887_1135 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1136 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h470 == _T_481) begin
          _T_6887_1136 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1137 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h471 == _T_481) begin
          _T_6887_1137 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1138 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h472 == _T_481) begin
          _T_6887_1138 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1139 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h473 == _T_481) begin
          _T_6887_1139 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1140 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h474 == _T_481) begin
          _T_6887_1140 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1141 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h475 == _T_481) begin
          _T_6887_1141 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1142 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h476 == _T_481) begin
          _T_6887_1142 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1143 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h477 == _T_481) begin
          _T_6887_1143 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1144 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h478 == _T_481) begin
          _T_6887_1144 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1145 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h479 == _T_481) begin
          _T_6887_1145 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1146 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47a == _T_481) begin
          _T_6887_1146 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1147 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47b == _T_481) begin
          _T_6887_1147 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1148 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47c == _T_481) begin
          _T_6887_1148 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1149 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47d == _T_481) begin
          _T_6887_1149 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1150 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47e == _T_481) begin
          _T_6887_1150 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1151 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h47f == _T_481) begin
          _T_6887_1151 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1152 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h480 == _T_481) begin
          _T_6887_1152 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1153 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h481 == _T_481) begin
          _T_6887_1153 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1154 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h482 == _T_481) begin
          _T_6887_1154 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1155 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h483 == _T_481) begin
          _T_6887_1155 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1156 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h484 == _T_481) begin
          _T_6887_1156 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1157 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h485 == _T_481) begin
          _T_6887_1157 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1158 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h486 == _T_481) begin
          _T_6887_1158 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1159 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h487 == _T_481) begin
          _T_6887_1159 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1160 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h488 == _T_481) begin
          _T_6887_1160 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1161 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h489 == _T_481) begin
          _T_6887_1161 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1162 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48a == _T_481) begin
          _T_6887_1162 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1163 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48b == _T_481) begin
          _T_6887_1163 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1164 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48c == _T_481) begin
          _T_6887_1164 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1165 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48d == _T_481) begin
          _T_6887_1165 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1166 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48e == _T_481) begin
          _T_6887_1166 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1167 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h48f == _T_481) begin
          _T_6887_1167 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1168 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h490 == _T_481) begin
          _T_6887_1168 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1169 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h491 == _T_481) begin
          _T_6887_1169 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1170 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h492 == _T_481) begin
          _T_6887_1170 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1171 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h493 == _T_481) begin
          _T_6887_1171 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1172 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h494 == _T_481) begin
          _T_6887_1172 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1173 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h495 == _T_481) begin
          _T_6887_1173 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1174 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h496 == _T_481) begin
          _T_6887_1174 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1175 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h497 == _T_481) begin
          _T_6887_1175 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1176 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h498 == _T_481) begin
          _T_6887_1176 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1177 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h499 == _T_481) begin
          _T_6887_1177 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1178 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49a == _T_481) begin
          _T_6887_1178 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1179 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49b == _T_481) begin
          _T_6887_1179 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1180 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49c == _T_481) begin
          _T_6887_1180 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1181 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49d == _T_481) begin
          _T_6887_1181 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1182 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49e == _T_481) begin
          _T_6887_1182 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1183 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h49f == _T_481) begin
          _T_6887_1183 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1184 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a0 == _T_481) begin
          _T_6887_1184 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1185 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a1 == _T_481) begin
          _T_6887_1185 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1186 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a2 == _T_481) begin
          _T_6887_1186 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1187 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a3 == _T_481) begin
          _T_6887_1187 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1188 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a4 == _T_481) begin
          _T_6887_1188 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1189 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a5 == _T_481) begin
          _T_6887_1189 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1190 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a6 == _T_481) begin
          _T_6887_1190 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1191 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a7 == _T_481) begin
          _T_6887_1191 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1192 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a8 == _T_481) begin
          _T_6887_1192 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1193 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4a9 == _T_481) begin
          _T_6887_1193 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1194 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4aa == _T_481) begin
          _T_6887_1194 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1195 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ab == _T_481) begin
          _T_6887_1195 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1196 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ac == _T_481) begin
          _T_6887_1196 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1197 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ad == _T_481) begin
          _T_6887_1197 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1198 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ae == _T_481) begin
          _T_6887_1198 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1199 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4af == _T_481) begin
          _T_6887_1199 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1200 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b0 == _T_481) begin
          _T_6887_1200 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1201 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b1 == _T_481) begin
          _T_6887_1201 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1202 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b2 == _T_481) begin
          _T_6887_1202 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1203 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b3 == _T_481) begin
          _T_6887_1203 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1204 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b4 == _T_481) begin
          _T_6887_1204 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1205 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b5 == _T_481) begin
          _T_6887_1205 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1206 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b6 == _T_481) begin
          _T_6887_1206 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1207 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b7 == _T_481) begin
          _T_6887_1207 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1208 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b8 == _T_481) begin
          _T_6887_1208 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1209 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4b9 == _T_481) begin
          _T_6887_1209 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1210 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ba == _T_481) begin
          _T_6887_1210 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1211 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4bb == _T_481) begin
          _T_6887_1211 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1212 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4bc == _T_481) begin
          _T_6887_1212 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1213 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4bd == _T_481) begin
          _T_6887_1213 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1214 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4be == _T_481) begin
          _T_6887_1214 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1215 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4bf == _T_481) begin
          _T_6887_1215 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1216 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c0 == _T_481) begin
          _T_6887_1216 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1217 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c1 == _T_481) begin
          _T_6887_1217 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1218 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c2 == _T_481) begin
          _T_6887_1218 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1219 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c3 == _T_481) begin
          _T_6887_1219 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1220 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c4 == _T_481) begin
          _T_6887_1220 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1221 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c5 == _T_481) begin
          _T_6887_1221 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1222 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c6 == _T_481) begin
          _T_6887_1222 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1223 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c7 == _T_481) begin
          _T_6887_1223 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1224 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c8 == _T_481) begin
          _T_6887_1224 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1225 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4c9 == _T_481) begin
          _T_6887_1225 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1226 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ca == _T_481) begin
          _T_6887_1226 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1227 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4cb == _T_481) begin
          _T_6887_1227 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1228 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4cc == _T_481) begin
          _T_6887_1228 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1229 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4cd == _T_481) begin
          _T_6887_1229 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1230 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ce == _T_481) begin
          _T_6887_1230 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1231 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4cf == _T_481) begin
          _T_6887_1231 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1232 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d0 == _T_481) begin
          _T_6887_1232 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1233 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d1 == _T_481) begin
          _T_6887_1233 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1234 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d2 == _T_481) begin
          _T_6887_1234 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1235 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d3 == _T_481) begin
          _T_6887_1235 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1236 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d4 == _T_481) begin
          _T_6887_1236 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1237 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d5 == _T_481) begin
          _T_6887_1237 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1238 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d6 == _T_481) begin
          _T_6887_1238 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1239 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d7 == _T_481) begin
          _T_6887_1239 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1240 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d8 == _T_481) begin
          _T_6887_1240 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1241 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4d9 == _T_481) begin
          _T_6887_1241 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1242 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4da == _T_481) begin
          _T_6887_1242 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1243 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4db == _T_481) begin
          _T_6887_1243 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1244 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4dc == _T_481) begin
          _T_6887_1244 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1245 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4dd == _T_481) begin
          _T_6887_1245 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1246 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4de == _T_481) begin
          _T_6887_1246 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1247 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4df == _T_481) begin
          _T_6887_1247 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1248 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e0 == _T_481) begin
          _T_6887_1248 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1249 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e1 == _T_481) begin
          _T_6887_1249 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1250 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e2 == _T_481) begin
          _T_6887_1250 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1251 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e3 == _T_481) begin
          _T_6887_1251 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1252 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e4 == _T_481) begin
          _T_6887_1252 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1253 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e5 == _T_481) begin
          _T_6887_1253 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1254 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e6 == _T_481) begin
          _T_6887_1254 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1255 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e7 == _T_481) begin
          _T_6887_1255 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1256 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e8 == _T_481) begin
          _T_6887_1256 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1257 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4e9 == _T_481) begin
          _T_6887_1257 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1258 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ea == _T_481) begin
          _T_6887_1258 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1259 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4eb == _T_481) begin
          _T_6887_1259 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1260 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ec == _T_481) begin
          _T_6887_1260 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1261 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ed == _T_481) begin
          _T_6887_1261 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1262 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ee == _T_481) begin
          _T_6887_1262 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1263 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ef == _T_481) begin
          _T_6887_1263 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1264 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f0 == _T_481) begin
          _T_6887_1264 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1265 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f1 == _T_481) begin
          _T_6887_1265 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1266 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f2 == _T_481) begin
          _T_6887_1266 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1267 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f3 == _T_481) begin
          _T_6887_1267 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1268 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f4 == _T_481) begin
          _T_6887_1268 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1269 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f5 == _T_481) begin
          _T_6887_1269 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1270 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f6 == _T_481) begin
          _T_6887_1270 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1271 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f7 == _T_481) begin
          _T_6887_1271 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1272 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f8 == _T_481) begin
          _T_6887_1272 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1273 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4f9 == _T_481) begin
          _T_6887_1273 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1274 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4fa == _T_481) begin
          _T_6887_1274 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1275 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4fb == _T_481) begin
          _T_6887_1275 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1276 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4fc == _T_481) begin
          _T_6887_1276 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1277 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4fd == _T_481) begin
          _T_6887_1277 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1278 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4fe == _T_481) begin
          _T_6887_1278 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1279 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h4ff == _T_481) begin
          _T_6887_1279 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1280 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h500 == _T_481) begin
          _T_6887_1280 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1281 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h501 == _T_481) begin
          _T_6887_1281 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1282 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h502 == _T_481) begin
          _T_6887_1282 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1283 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h503 == _T_481) begin
          _T_6887_1283 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1284 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h504 == _T_481) begin
          _T_6887_1284 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1285 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h505 == _T_481) begin
          _T_6887_1285 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1286 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h506 == _T_481) begin
          _T_6887_1286 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1287 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h507 == _T_481) begin
          _T_6887_1287 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1288 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h508 == _T_481) begin
          _T_6887_1288 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1289 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h509 == _T_481) begin
          _T_6887_1289 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1290 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50a == _T_481) begin
          _T_6887_1290 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1291 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50b == _T_481) begin
          _T_6887_1291 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1292 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50c == _T_481) begin
          _T_6887_1292 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1293 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50d == _T_481) begin
          _T_6887_1293 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1294 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50e == _T_481) begin
          _T_6887_1294 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1295 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h50f == _T_481) begin
          _T_6887_1295 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1296 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h510 == _T_481) begin
          _T_6887_1296 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1297 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h511 == _T_481) begin
          _T_6887_1297 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1298 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h512 == _T_481) begin
          _T_6887_1298 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1299 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h513 == _T_481) begin
          _T_6887_1299 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1300 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h514 == _T_481) begin
          _T_6887_1300 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1301 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h515 == _T_481) begin
          _T_6887_1301 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1302 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h516 == _T_481) begin
          _T_6887_1302 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1303 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h517 == _T_481) begin
          _T_6887_1303 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1304 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h518 == _T_481) begin
          _T_6887_1304 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1305 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h519 == _T_481) begin
          _T_6887_1305 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1306 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51a == _T_481) begin
          _T_6887_1306 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1307 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51b == _T_481) begin
          _T_6887_1307 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1308 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51c == _T_481) begin
          _T_6887_1308 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1309 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51d == _T_481) begin
          _T_6887_1309 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1310 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51e == _T_481) begin
          _T_6887_1310 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1311 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h51f == _T_481) begin
          _T_6887_1311 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1312 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h520 == _T_481) begin
          _T_6887_1312 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1313 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h521 == _T_481) begin
          _T_6887_1313 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1314 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h522 == _T_481) begin
          _T_6887_1314 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1315 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h523 == _T_481) begin
          _T_6887_1315 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1316 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h524 == _T_481) begin
          _T_6887_1316 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1317 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h525 == _T_481) begin
          _T_6887_1317 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1318 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h526 == _T_481) begin
          _T_6887_1318 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1319 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h527 == _T_481) begin
          _T_6887_1319 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1320 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h528 == _T_481) begin
          _T_6887_1320 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1321 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h529 == _T_481) begin
          _T_6887_1321 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1322 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52a == _T_481) begin
          _T_6887_1322 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1323 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52b == _T_481) begin
          _T_6887_1323 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1324 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52c == _T_481) begin
          _T_6887_1324 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1325 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52d == _T_481) begin
          _T_6887_1325 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1326 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52e == _T_481) begin
          _T_6887_1326 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1327 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h52f == _T_481) begin
          _T_6887_1327 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1328 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h530 == _T_481) begin
          _T_6887_1328 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1329 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h531 == _T_481) begin
          _T_6887_1329 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1330 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h532 == _T_481) begin
          _T_6887_1330 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1331 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h533 == _T_481) begin
          _T_6887_1331 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1332 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h534 == _T_481) begin
          _T_6887_1332 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1333 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h535 == _T_481) begin
          _T_6887_1333 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1334 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h536 == _T_481) begin
          _T_6887_1334 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1335 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h537 == _T_481) begin
          _T_6887_1335 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1336 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h538 == _T_481) begin
          _T_6887_1336 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1337 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h539 == _T_481) begin
          _T_6887_1337 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1338 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53a == _T_481) begin
          _T_6887_1338 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1339 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53b == _T_481) begin
          _T_6887_1339 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1340 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53c == _T_481) begin
          _T_6887_1340 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1341 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53d == _T_481) begin
          _T_6887_1341 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1342 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53e == _T_481) begin
          _T_6887_1342 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1343 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h53f == _T_481) begin
          _T_6887_1343 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1344 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h540 == _T_481) begin
          _T_6887_1344 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1345 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h541 == _T_481) begin
          _T_6887_1345 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1346 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h542 == _T_481) begin
          _T_6887_1346 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1347 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h543 == _T_481) begin
          _T_6887_1347 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1348 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h544 == _T_481) begin
          _T_6887_1348 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1349 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h545 == _T_481) begin
          _T_6887_1349 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1350 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h546 == _T_481) begin
          _T_6887_1350 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1351 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h547 == _T_481) begin
          _T_6887_1351 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1352 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h548 == _T_481) begin
          _T_6887_1352 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1353 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h549 == _T_481) begin
          _T_6887_1353 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1354 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54a == _T_481) begin
          _T_6887_1354 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1355 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54b == _T_481) begin
          _T_6887_1355 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1356 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54c == _T_481) begin
          _T_6887_1356 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1357 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54d == _T_481) begin
          _T_6887_1357 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1358 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54e == _T_481) begin
          _T_6887_1358 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1359 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h54f == _T_481) begin
          _T_6887_1359 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1360 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h550 == _T_481) begin
          _T_6887_1360 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1361 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h551 == _T_481) begin
          _T_6887_1361 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1362 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h552 == _T_481) begin
          _T_6887_1362 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1363 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h553 == _T_481) begin
          _T_6887_1363 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1364 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h554 == _T_481) begin
          _T_6887_1364 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1365 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h555 == _T_481) begin
          _T_6887_1365 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1366 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h556 == _T_481) begin
          _T_6887_1366 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1367 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h557 == _T_481) begin
          _T_6887_1367 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1368 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h558 == _T_481) begin
          _T_6887_1368 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1369 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h559 == _T_481) begin
          _T_6887_1369 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1370 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55a == _T_481) begin
          _T_6887_1370 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1371 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55b == _T_481) begin
          _T_6887_1371 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1372 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55c == _T_481) begin
          _T_6887_1372 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1373 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55d == _T_481) begin
          _T_6887_1373 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1374 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55e == _T_481) begin
          _T_6887_1374 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1375 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h55f == _T_481) begin
          _T_6887_1375 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1376 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h560 == _T_481) begin
          _T_6887_1376 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1377 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h561 == _T_481) begin
          _T_6887_1377 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1378 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h562 == _T_481) begin
          _T_6887_1378 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1379 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h563 == _T_481) begin
          _T_6887_1379 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1380 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h564 == _T_481) begin
          _T_6887_1380 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1381 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h565 == _T_481) begin
          _T_6887_1381 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1382 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h566 == _T_481) begin
          _T_6887_1382 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1383 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h567 == _T_481) begin
          _T_6887_1383 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1384 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h568 == _T_481) begin
          _T_6887_1384 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1385 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h569 == _T_481) begin
          _T_6887_1385 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1386 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56a == _T_481) begin
          _T_6887_1386 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1387 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56b == _T_481) begin
          _T_6887_1387 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1388 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56c == _T_481) begin
          _T_6887_1388 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1389 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56d == _T_481) begin
          _T_6887_1389 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1390 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56e == _T_481) begin
          _T_6887_1390 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1391 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h56f == _T_481) begin
          _T_6887_1391 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1392 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h570 == _T_481) begin
          _T_6887_1392 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1393 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h571 == _T_481) begin
          _T_6887_1393 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1394 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h572 == _T_481) begin
          _T_6887_1394 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1395 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h573 == _T_481) begin
          _T_6887_1395 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1396 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h574 == _T_481) begin
          _T_6887_1396 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1397 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h575 == _T_481) begin
          _T_6887_1397 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1398 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h576 == _T_481) begin
          _T_6887_1398 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1399 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h577 == _T_481) begin
          _T_6887_1399 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1400 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h578 == _T_481) begin
          _T_6887_1400 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1401 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h579 == _T_481) begin
          _T_6887_1401 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1402 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57a == _T_481) begin
          _T_6887_1402 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1403 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57b == _T_481) begin
          _T_6887_1403 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1404 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57c == _T_481) begin
          _T_6887_1404 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1405 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57d == _T_481) begin
          _T_6887_1405 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1406 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57e == _T_481) begin
          _T_6887_1406 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1407 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h57f == _T_481) begin
          _T_6887_1407 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1408 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h580 == _T_481) begin
          _T_6887_1408 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1409 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h581 == _T_481) begin
          _T_6887_1409 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1410 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h582 == _T_481) begin
          _T_6887_1410 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1411 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h583 == _T_481) begin
          _T_6887_1411 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1412 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h584 == _T_481) begin
          _T_6887_1412 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1413 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h585 == _T_481) begin
          _T_6887_1413 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1414 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h586 == _T_481) begin
          _T_6887_1414 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1415 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h587 == _T_481) begin
          _T_6887_1415 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1416 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h588 == _T_481) begin
          _T_6887_1416 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1417 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h589 == _T_481) begin
          _T_6887_1417 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1418 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58a == _T_481) begin
          _T_6887_1418 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1419 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58b == _T_481) begin
          _T_6887_1419 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1420 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58c == _T_481) begin
          _T_6887_1420 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1421 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58d == _T_481) begin
          _T_6887_1421 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1422 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58e == _T_481) begin
          _T_6887_1422 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1423 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h58f == _T_481) begin
          _T_6887_1423 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1424 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h590 == _T_481) begin
          _T_6887_1424 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1425 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h591 == _T_481) begin
          _T_6887_1425 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1426 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h592 == _T_481) begin
          _T_6887_1426 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1427 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h593 == _T_481) begin
          _T_6887_1427 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1428 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h594 == _T_481) begin
          _T_6887_1428 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1429 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h595 == _T_481) begin
          _T_6887_1429 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1430 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h596 == _T_481) begin
          _T_6887_1430 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1431 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h597 == _T_481) begin
          _T_6887_1431 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1432 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h598 == _T_481) begin
          _T_6887_1432 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1433 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h599 == _T_481) begin
          _T_6887_1433 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1434 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59a == _T_481) begin
          _T_6887_1434 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1435 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59b == _T_481) begin
          _T_6887_1435 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1436 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59c == _T_481) begin
          _T_6887_1436 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1437 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59d == _T_481) begin
          _T_6887_1437 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1438 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59e == _T_481) begin
          _T_6887_1438 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1439 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h59f == _T_481) begin
          _T_6887_1439 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1440 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a0 == _T_481) begin
          _T_6887_1440 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1441 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a1 == _T_481) begin
          _T_6887_1441 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1442 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a2 == _T_481) begin
          _T_6887_1442 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1443 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a3 == _T_481) begin
          _T_6887_1443 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1444 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a4 == _T_481) begin
          _T_6887_1444 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1445 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a5 == _T_481) begin
          _T_6887_1445 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1446 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a6 == _T_481) begin
          _T_6887_1446 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1447 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a7 == _T_481) begin
          _T_6887_1447 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1448 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a8 == _T_481) begin
          _T_6887_1448 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1449 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5a9 == _T_481) begin
          _T_6887_1449 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1450 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5aa == _T_481) begin
          _T_6887_1450 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1451 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ab == _T_481) begin
          _T_6887_1451 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1452 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ac == _T_481) begin
          _T_6887_1452 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1453 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ad == _T_481) begin
          _T_6887_1453 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1454 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ae == _T_481) begin
          _T_6887_1454 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1455 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5af == _T_481) begin
          _T_6887_1455 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1456 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b0 == _T_481) begin
          _T_6887_1456 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1457 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b1 == _T_481) begin
          _T_6887_1457 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1458 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b2 == _T_481) begin
          _T_6887_1458 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1459 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b3 == _T_481) begin
          _T_6887_1459 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1460 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b4 == _T_481) begin
          _T_6887_1460 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1461 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b5 == _T_481) begin
          _T_6887_1461 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1462 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b6 == _T_481) begin
          _T_6887_1462 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1463 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b7 == _T_481) begin
          _T_6887_1463 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1464 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b8 == _T_481) begin
          _T_6887_1464 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1465 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5b9 == _T_481) begin
          _T_6887_1465 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1466 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ba == _T_481) begin
          _T_6887_1466 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1467 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5bb == _T_481) begin
          _T_6887_1467 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1468 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5bc == _T_481) begin
          _T_6887_1468 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1469 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5bd == _T_481) begin
          _T_6887_1469 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1470 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5be == _T_481) begin
          _T_6887_1470 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1471 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5bf == _T_481) begin
          _T_6887_1471 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1472 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c0 == _T_481) begin
          _T_6887_1472 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1473 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c1 == _T_481) begin
          _T_6887_1473 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1474 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c2 == _T_481) begin
          _T_6887_1474 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1475 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c3 == _T_481) begin
          _T_6887_1475 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1476 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c4 == _T_481) begin
          _T_6887_1476 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1477 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c5 == _T_481) begin
          _T_6887_1477 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1478 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c6 == _T_481) begin
          _T_6887_1478 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1479 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c7 == _T_481) begin
          _T_6887_1479 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1480 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c8 == _T_481) begin
          _T_6887_1480 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1481 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5c9 == _T_481) begin
          _T_6887_1481 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1482 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ca == _T_481) begin
          _T_6887_1482 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1483 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5cb == _T_481) begin
          _T_6887_1483 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1484 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5cc == _T_481) begin
          _T_6887_1484 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1485 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5cd == _T_481) begin
          _T_6887_1485 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1486 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ce == _T_481) begin
          _T_6887_1486 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1487 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5cf == _T_481) begin
          _T_6887_1487 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1488 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d0 == _T_481) begin
          _T_6887_1488 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1489 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d1 == _T_481) begin
          _T_6887_1489 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1490 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d2 == _T_481) begin
          _T_6887_1490 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1491 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d3 == _T_481) begin
          _T_6887_1491 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1492 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d4 == _T_481) begin
          _T_6887_1492 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1493 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d5 == _T_481) begin
          _T_6887_1493 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1494 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d6 == _T_481) begin
          _T_6887_1494 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1495 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d7 == _T_481) begin
          _T_6887_1495 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1496 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d8 == _T_481) begin
          _T_6887_1496 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1497 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5d9 == _T_481) begin
          _T_6887_1497 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1498 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5da == _T_481) begin
          _T_6887_1498 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1499 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5db == _T_481) begin
          _T_6887_1499 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1500 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5dc == _T_481) begin
          _T_6887_1500 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1501 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5dd == _T_481) begin
          _T_6887_1501 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1502 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5de == _T_481) begin
          _T_6887_1502 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1503 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5df == _T_481) begin
          _T_6887_1503 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1504 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e0 == _T_481) begin
          _T_6887_1504 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1505 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e1 == _T_481) begin
          _T_6887_1505 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1506 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e2 == _T_481) begin
          _T_6887_1506 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1507 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e3 == _T_481) begin
          _T_6887_1507 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1508 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e4 == _T_481) begin
          _T_6887_1508 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1509 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e5 == _T_481) begin
          _T_6887_1509 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1510 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e6 == _T_481) begin
          _T_6887_1510 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1511 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e7 == _T_481) begin
          _T_6887_1511 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1512 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e8 == _T_481) begin
          _T_6887_1512 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1513 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5e9 == _T_481) begin
          _T_6887_1513 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1514 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ea == _T_481) begin
          _T_6887_1514 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1515 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5eb == _T_481) begin
          _T_6887_1515 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1516 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ec == _T_481) begin
          _T_6887_1516 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1517 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ed == _T_481) begin
          _T_6887_1517 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1518 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ee == _T_481) begin
          _T_6887_1518 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1519 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ef == _T_481) begin
          _T_6887_1519 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1520 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f0 == _T_481) begin
          _T_6887_1520 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1521 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f1 == _T_481) begin
          _T_6887_1521 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1522 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f2 == _T_481) begin
          _T_6887_1522 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1523 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f3 == _T_481) begin
          _T_6887_1523 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1524 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f4 == _T_481) begin
          _T_6887_1524 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1525 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f5 == _T_481) begin
          _T_6887_1525 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1526 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f6 == _T_481) begin
          _T_6887_1526 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1527 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f7 == _T_481) begin
          _T_6887_1527 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1528 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f8 == _T_481) begin
          _T_6887_1528 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1529 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5f9 == _T_481) begin
          _T_6887_1529 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1530 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5fa == _T_481) begin
          _T_6887_1530 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1531 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5fb == _T_481) begin
          _T_6887_1531 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1532 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5fc == _T_481) begin
          _T_6887_1532 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1533 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5fd == _T_481) begin
          _T_6887_1533 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1534 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5fe == _T_481) begin
          _T_6887_1534 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1535 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h5ff == _T_481) begin
          _T_6887_1535 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1536 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h600 == _T_481) begin
          _T_6887_1536 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1537 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h601 == _T_481) begin
          _T_6887_1537 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1538 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h602 == _T_481) begin
          _T_6887_1538 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1539 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h603 == _T_481) begin
          _T_6887_1539 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1540 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h604 == _T_481) begin
          _T_6887_1540 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1541 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h605 == _T_481) begin
          _T_6887_1541 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1542 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h606 == _T_481) begin
          _T_6887_1542 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1543 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h607 == _T_481) begin
          _T_6887_1543 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1544 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h608 == _T_481) begin
          _T_6887_1544 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1545 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h609 == _T_481) begin
          _T_6887_1545 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1546 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60a == _T_481) begin
          _T_6887_1546 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1547 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60b == _T_481) begin
          _T_6887_1547 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1548 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60c == _T_481) begin
          _T_6887_1548 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1549 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60d == _T_481) begin
          _T_6887_1549 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1550 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60e == _T_481) begin
          _T_6887_1550 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1551 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h60f == _T_481) begin
          _T_6887_1551 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1552 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h610 == _T_481) begin
          _T_6887_1552 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1553 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h611 == _T_481) begin
          _T_6887_1553 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1554 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h612 == _T_481) begin
          _T_6887_1554 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1555 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h613 == _T_481) begin
          _T_6887_1555 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1556 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h614 == _T_481) begin
          _T_6887_1556 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1557 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h615 == _T_481) begin
          _T_6887_1557 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1558 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h616 == _T_481) begin
          _T_6887_1558 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1559 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h617 == _T_481) begin
          _T_6887_1559 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1560 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h618 == _T_481) begin
          _T_6887_1560 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1561 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h619 == _T_481) begin
          _T_6887_1561 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1562 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61a == _T_481) begin
          _T_6887_1562 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1563 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61b == _T_481) begin
          _T_6887_1563 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1564 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61c == _T_481) begin
          _T_6887_1564 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1565 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61d == _T_481) begin
          _T_6887_1565 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1566 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61e == _T_481) begin
          _T_6887_1566 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1567 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h61f == _T_481) begin
          _T_6887_1567 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1568 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h620 == _T_481) begin
          _T_6887_1568 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1569 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h621 == _T_481) begin
          _T_6887_1569 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1570 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h622 == _T_481) begin
          _T_6887_1570 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1571 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h623 == _T_481) begin
          _T_6887_1571 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1572 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h624 == _T_481) begin
          _T_6887_1572 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1573 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h625 == _T_481) begin
          _T_6887_1573 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1574 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h626 == _T_481) begin
          _T_6887_1574 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1575 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h627 == _T_481) begin
          _T_6887_1575 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1576 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h628 == _T_481) begin
          _T_6887_1576 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1577 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h629 == _T_481) begin
          _T_6887_1577 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1578 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62a == _T_481) begin
          _T_6887_1578 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1579 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62b == _T_481) begin
          _T_6887_1579 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1580 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62c == _T_481) begin
          _T_6887_1580 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1581 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62d == _T_481) begin
          _T_6887_1581 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1582 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62e == _T_481) begin
          _T_6887_1582 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1583 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h62f == _T_481) begin
          _T_6887_1583 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1584 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h630 == _T_481) begin
          _T_6887_1584 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1585 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h631 == _T_481) begin
          _T_6887_1585 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1586 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h632 == _T_481) begin
          _T_6887_1586 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1587 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h633 == _T_481) begin
          _T_6887_1587 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1588 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h634 == _T_481) begin
          _T_6887_1588 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1589 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h635 == _T_481) begin
          _T_6887_1589 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1590 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h636 == _T_481) begin
          _T_6887_1590 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1591 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h637 == _T_481) begin
          _T_6887_1591 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1592 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h638 == _T_481) begin
          _T_6887_1592 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1593 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h639 == _T_481) begin
          _T_6887_1593 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1594 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63a == _T_481) begin
          _T_6887_1594 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1595 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63b == _T_481) begin
          _T_6887_1595 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1596 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63c == _T_481) begin
          _T_6887_1596 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1597 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63d == _T_481) begin
          _T_6887_1597 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1598 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63e == _T_481) begin
          _T_6887_1598 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1599 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h63f == _T_481) begin
          _T_6887_1599 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1600 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h640 == _T_481) begin
          _T_6887_1600 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1601 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h641 == _T_481) begin
          _T_6887_1601 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1602 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h642 == _T_481) begin
          _T_6887_1602 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1603 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h643 == _T_481) begin
          _T_6887_1603 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1604 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h644 == _T_481) begin
          _T_6887_1604 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1605 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h645 == _T_481) begin
          _T_6887_1605 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1606 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h646 == _T_481) begin
          _T_6887_1606 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1607 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h647 == _T_481) begin
          _T_6887_1607 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1608 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h648 == _T_481) begin
          _T_6887_1608 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1609 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h649 == _T_481) begin
          _T_6887_1609 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1610 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64a == _T_481) begin
          _T_6887_1610 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1611 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64b == _T_481) begin
          _T_6887_1611 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1612 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64c == _T_481) begin
          _T_6887_1612 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1613 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64d == _T_481) begin
          _T_6887_1613 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1614 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64e == _T_481) begin
          _T_6887_1614 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1615 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h64f == _T_481) begin
          _T_6887_1615 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1616 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h650 == _T_481) begin
          _T_6887_1616 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1617 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h651 == _T_481) begin
          _T_6887_1617 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1618 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h652 == _T_481) begin
          _T_6887_1618 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1619 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h653 == _T_481) begin
          _T_6887_1619 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1620 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h654 == _T_481) begin
          _T_6887_1620 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1621 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h655 == _T_481) begin
          _T_6887_1621 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1622 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h656 == _T_481) begin
          _T_6887_1622 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1623 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h657 == _T_481) begin
          _T_6887_1623 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1624 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h658 == _T_481) begin
          _T_6887_1624 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1625 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h659 == _T_481) begin
          _T_6887_1625 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1626 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65a == _T_481) begin
          _T_6887_1626 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1627 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65b == _T_481) begin
          _T_6887_1627 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1628 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65c == _T_481) begin
          _T_6887_1628 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1629 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65d == _T_481) begin
          _T_6887_1629 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1630 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65e == _T_481) begin
          _T_6887_1630 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1631 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h65f == _T_481) begin
          _T_6887_1631 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1632 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h660 == _T_481) begin
          _T_6887_1632 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1633 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h661 == _T_481) begin
          _T_6887_1633 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1634 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h662 == _T_481) begin
          _T_6887_1634 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1635 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h663 == _T_481) begin
          _T_6887_1635 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1636 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h664 == _T_481) begin
          _T_6887_1636 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1637 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h665 == _T_481) begin
          _T_6887_1637 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1638 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h666 == _T_481) begin
          _T_6887_1638 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1639 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h667 == _T_481) begin
          _T_6887_1639 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1640 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h668 == _T_481) begin
          _T_6887_1640 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1641 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h669 == _T_481) begin
          _T_6887_1641 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1642 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66a == _T_481) begin
          _T_6887_1642 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1643 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66b == _T_481) begin
          _T_6887_1643 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1644 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66c == _T_481) begin
          _T_6887_1644 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1645 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66d == _T_481) begin
          _T_6887_1645 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1646 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66e == _T_481) begin
          _T_6887_1646 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1647 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h66f == _T_481) begin
          _T_6887_1647 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1648 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h670 == _T_481) begin
          _T_6887_1648 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1649 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h671 == _T_481) begin
          _T_6887_1649 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1650 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h672 == _T_481) begin
          _T_6887_1650 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1651 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h673 == _T_481) begin
          _T_6887_1651 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1652 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h674 == _T_481) begin
          _T_6887_1652 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1653 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h675 == _T_481) begin
          _T_6887_1653 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1654 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h676 == _T_481) begin
          _T_6887_1654 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1655 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h677 == _T_481) begin
          _T_6887_1655 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1656 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h678 == _T_481) begin
          _T_6887_1656 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1657 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h679 == _T_481) begin
          _T_6887_1657 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1658 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67a == _T_481) begin
          _T_6887_1658 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1659 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67b == _T_481) begin
          _T_6887_1659 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1660 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67c == _T_481) begin
          _T_6887_1660 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1661 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67d == _T_481) begin
          _T_6887_1661 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1662 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67e == _T_481) begin
          _T_6887_1662 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1663 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h67f == _T_481) begin
          _T_6887_1663 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1664 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h680 == _T_481) begin
          _T_6887_1664 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1665 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h681 == _T_481) begin
          _T_6887_1665 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1666 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h682 == _T_481) begin
          _T_6887_1666 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1667 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h683 == _T_481) begin
          _T_6887_1667 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1668 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h684 == _T_481) begin
          _T_6887_1668 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1669 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h685 == _T_481) begin
          _T_6887_1669 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1670 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h686 == _T_481) begin
          _T_6887_1670 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1671 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h687 == _T_481) begin
          _T_6887_1671 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1672 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h688 == _T_481) begin
          _T_6887_1672 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1673 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h689 == _T_481) begin
          _T_6887_1673 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1674 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68a == _T_481) begin
          _T_6887_1674 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1675 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68b == _T_481) begin
          _T_6887_1675 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1676 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68c == _T_481) begin
          _T_6887_1676 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1677 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68d == _T_481) begin
          _T_6887_1677 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1678 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68e == _T_481) begin
          _T_6887_1678 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1679 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h68f == _T_481) begin
          _T_6887_1679 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1680 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h690 == _T_481) begin
          _T_6887_1680 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1681 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h691 == _T_481) begin
          _T_6887_1681 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1682 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h692 == _T_481) begin
          _T_6887_1682 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1683 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h693 == _T_481) begin
          _T_6887_1683 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1684 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h694 == _T_481) begin
          _T_6887_1684 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1685 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h695 == _T_481) begin
          _T_6887_1685 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1686 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h696 == _T_481) begin
          _T_6887_1686 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1687 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h697 == _T_481) begin
          _T_6887_1687 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1688 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h698 == _T_481) begin
          _T_6887_1688 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1689 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h699 == _T_481) begin
          _T_6887_1689 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1690 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69a == _T_481) begin
          _T_6887_1690 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1691 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69b == _T_481) begin
          _T_6887_1691 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1692 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69c == _T_481) begin
          _T_6887_1692 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1693 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69d == _T_481) begin
          _T_6887_1693 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1694 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69e == _T_481) begin
          _T_6887_1694 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1695 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h69f == _T_481) begin
          _T_6887_1695 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1696 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a0 == _T_481) begin
          _T_6887_1696 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1697 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a1 == _T_481) begin
          _T_6887_1697 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1698 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a2 == _T_481) begin
          _T_6887_1698 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1699 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a3 == _T_481) begin
          _T_6887_1699 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1700 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a4 == _T_481) begin
          _T_6887_1700 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1701 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a5 == _T_481) begin
          _T_6887_1701 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1702 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a6 == _T_481) begin
          _T_6887_1702 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1703 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a7 == _T_481) begin
          _T_6887_1703 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1704 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a8 == _T_481) begin
          _T_6887_1704 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1705 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6a9 == _T_481) begin
          _T_6887_1705 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1706 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6aa == _T_481) begin
          _T_6887_1706 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1707 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ab == _T_481) begin
          _T_6887_1707 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1708 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ac == _T_481) begin
          _T_6887_1708 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1709 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ad == _T_481) begin
          _T_6887_1709 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1710 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ae == _T_481) begin
          _T_6887_1710 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1711 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6af == _T_481) begin
          _T_6887_1711 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1712 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b0 == _T_481) begin
          _T_6887_1712 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1713 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b1 == _T_481) begin
          _T_6887_1713 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1714 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b2 == _T_481) begin
          _T_6887_1714 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1715 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b3 == _T_481) begin
          _T_6887_1715 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1716 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b4 == _T_481) begin
          _T_6887_1716 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1717 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b5 == _T_481) begin
          _T_6887_1717 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1718 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b6 == _T_481) begin
          _T_6887_1718 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1719 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b7 == _T_481) begin
          _T_6887_1719 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1720 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b8 == _T_481) begin
          _T_6887_1720 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1721 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6b9 == _T_481) begin
          _T_6887_1721 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1722 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ba == _T_481) begin
          _T_6887_1722 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1723 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6bb == _T_481) begin
          _T_6887_1723 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1724 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6bc == _T_481) begin
          _T_6887_1724 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1725 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6bd == _T_481) begin
          _T_6887_1725 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1726 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6be == _T_481) begin
          _T_6887_1726 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1727 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6bf == _T_481) begin
          _T_6887_1727 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1728 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c0 == _T_481) begin
          _T_6887_1728 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1729 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c1 == _T_481) begin
          _T_6887_1729 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1730 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c2 == _T_481) begin
          _T_6887_1730 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1731 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c3 == _T_481) begin
          _T_6887_1731 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1732 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c4 == _T_481) begin
          _T_6887_1732 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1733 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c5 == _T_481) begin
          _T_6887_1733 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1734 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c6 == _T_481) begin
          _T_6887_1734 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1735 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c7 == _T_481) begin
          _T_6887_1735 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1736 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c8 == _T_481) begin
          _T_6887_1736 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1737 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6c9 == _T_481) begin
          _T_6887_1737 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1738 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ca == _T_481) begin
          _T_6887_1738 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1739 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6cb == _T_481) begin
          _T_6887_1739 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1740 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6cc == _T_481) begin
          _T_6887_1740 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1741 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6cd == _T_481) begin
          _T_6887_1741 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1742 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ce == _T_481) begin
          _T_6887_1742 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1743 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6cf == _T_481) begin
          _T_6887_1743 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1744 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d0 == _T_481) begin
          _T_6887_1744 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1745 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d1 == _T_481) begin
          _T_6887_1745 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1746 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d2 == _T_481) begin
          _T_6887_1746 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1747 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d3 == _T_481) begin
          _T_6887_1747 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1748 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d4 == _T_481) begin
          _T_6887_1748 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1749 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d5 == _T_481) begin
          _T_6887_1749 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1750 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d6 == _T_481) begin
          _T_6887_1750 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1751 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d7 == _T_481) begin
          _T_6887_1751 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1752 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d8 == _T_481) begin
          _T_6887_1752 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1753 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6d9 == _T_481) begin
          _T_6887_1753 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1754 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6da == _T_481) begin
          _T_6887_1754 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1755 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6db == _T_481) begin
          _T_6887_1755 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1756 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6dc == _T_481) begin
          _T_6887_1756 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1757 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6dd == _T_481) begin
          _T_6887_1757 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1758 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6de == _T_481) begin
          _T_6887_1758 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1759 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6df == _T_481) begin
          _T_6887_1759 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1760 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e0 == _T_481) begin
          _T_6887_1760 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1761 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e1 == _T_481) begin
          _T_6887_1761 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1762 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e2 == _T_481) begin
          _T_6887_1762 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1763 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e3 == _T_481) begin
          _T_6887_1763 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1764 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e4 == _T_481) begin
          _T_6887_1764 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1765 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e5 == _T_481) begin
          _T_6887_1765 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1766 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e6 == _T_481) begin
          _T_6887_1766 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1767 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e7 == _T_481) begin
          _T_6887_1767 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1768 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e8 == _T_481) begin
          _T_6887_1768 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1769 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6e9 == _T_481) begin
          _T_6887_1769 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1770 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ea == _T_481) begin
          _T_6887_1770 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1771 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6eb == _T_481) begin
          _T_6887_1771 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1772 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ec == _T_481) begin
          _T_6887_1772 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1773 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ed == _T_481) begin
          _T_6887_1773 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1774 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ee == _T_481) begin
          _T_6887_1774 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1775 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ef == _T_481) begin
          _T_6887_1775 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1776 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f0 == _T_481) begin
          _T_6887_1776 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1777 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f1 == _T_481) begin
          _T_6887_1777 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1778 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f2 == _T_481) begin
          _T_6887_1778 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1779 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f3 == _T_481) begin
          _T_6887_1779 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1780 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f4 == _T_481) begin
          _T_6887_1780 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1781 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f5 == _T_481) begin
          _T_6887_1781 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1782 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f6 == _T_481) begin
          _T_6887_1782 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1783 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f7 == _T_481) begin
          _T_6887_1783 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1784 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f8 == _T_481) begin
          _T_6887_1784 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1785 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6f9 == _T_481) begin
          _T_6887_1785 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1786 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6fa == _T_481) begin
          _T_6887_1786 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1787 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6fb == _T_481) begin
          _T_6887_1787 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1788 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6fc == _T_481) begin
          _T_6887_1788 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1789 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6fd == _T_481) begin
          _T_6887_1789 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1790 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6fe == _T_481) begin
          _T_6887_1790 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1791 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h6ff == _T_481) begin
          _T_6887_1791 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1792 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h700 == _T_481) begin
          _T_6887_1792 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1793 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h701 == _T_481) begin
          _T_6887_1793 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1794 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h702 == _T_481) begin
          _T_6887_1794 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1795 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h703 == _T_481) begin
          _T_6887_1795 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1796 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h704 == _T_481) begin
          _T_6887_1796 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1797 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h705 == _T_481) begin
          _T_6887_1797 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1798 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h706 == _T_481) begin
          _T_6887_1798 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1799 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h707 == _T_481) begin
          _T_6887_1799 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1800 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h708 == _T_481) begin
          _T_6887_1800 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1801 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h709 == _T_481) begin
          _T_6887_1801 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1802 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70a == _T_481) begin
          _T_6887_1802 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1803 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70b == _T_481) begin
          _T_6887_1803 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1804 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70c == _T_481) begin
          _T_6887_1804 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1805 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70d == _T_481) begin
          _T_6887_1805 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1806 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70e == _T_481) begin
          _T_6887_1806 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1807 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h70f == _T_481) begin
          _T_6887_1807 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1808 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h710 == _T_481) begin
          _T_6887_1808 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1809 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h711 == _T_481) begin
          _T_6887_1809 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1810 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h712 == _T_481) begin
          _T_6887_1810 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1811 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h713 == _T_481) begin
          _T_6887_1811 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1812 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h714 == _T_481) begin
          _T_6887_1812 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1813 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h715 == _T_481) begin
          _T_6887_1813 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1814 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h716 == _T_481) begin
          _T_6887_1814 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1815 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h717 == _T_481) begin
          _T_6887_1815 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1816 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h718 == _T_481) begin
          _T_6887_1816 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1817 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h719 == _T_481) begin
          _T_6887_1817 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1818 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71a == _T_481) begin
          _T_6887_1818 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1819 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71b == _T_481) begin
          _T_6887_1819 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1820 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71c == _T_481) begin
          _T_6887_1820 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1821 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71d == _T_481) begin
          _T_6887_1821 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1822 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71e == _T_481) begin
          _T_6887_1822 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1823 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h71f == _T_481) begin
          _T_6887_1823 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1824 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h720 == _T_481) begin
          _T_6887_1824 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1825 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h721 == _T_481) begin
          _T_6887_1825 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1826 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h722 == _T_481) begin
          _T_6887_1826 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1827 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h723 == _T_481) begin
          _T_6887_1827 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1828 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h724 == _T_481) begin
          _T_6887_1828 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1829 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h725 == _T_481) begin
          _T_6887_1829 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1830 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h726 == _T_481) begin
          _T_6887_1830 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1831 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h727 == _T_481) begin
          _T_6887_1831 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1832 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h728 == _T_481) begin
          _T_6887_1832 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1833 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h729 == _T_481) begin
          _T_6887_1833 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1834 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72a == _T_481) begin
          _T_6887_1834 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1835 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72b == _T_481) begin
          _T_6887_1835 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1836 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72c == _T_481) begin
          _T_6887_1836 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1837 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72d == _T_481) begin
          _T_6887_1837 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1838 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72e == _T_481) begin
          _T_6887_1838 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1839 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h72f == _T_481) begin
          _T_6887_1839 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1840 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h730 == _T_481) begin
          _T_6887_1840 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1841 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h731 == _T_481) begin
          _T_6887_1841 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1842 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h732 == _T_481) begin
          _T_6887_1842 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1843 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h733 == _T_481) begin
          _T_6887_1843 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1844 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h734 == _T_481) begin
          _T_6887_1844 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1845 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h735 == _T_481) begin
          _T_6887_1845 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1846 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h736 == _T_481) begin
          _T_6887_1846 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1847 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h737 == _T_481) begin
          _T_6887_1847 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1848 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h738 == _T_481) begin
          _T_6887_1848 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1849 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h739 == _T_481) begin
          _T_6887_1849 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1850 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73a == _T_481) begin
          _T_6887_1850 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1851 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73b == _T_481) begin
          _T_6887_1851 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1852 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73c == _T_481) begin
          _T_6887_1852 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1853 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73d == _T_481) begin
          _T_6887_1853 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1854 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73e == _T_481) begin
          _T_6887_1854 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1855 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h73f == _T_481) begin
          _T_6887_1855 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1856 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h740 == _T_481) begin
          _T_6887_1856 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1857 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h741 == _T_481) begin
          _T_6887_1857 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1858 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h742 == _T_481) begin
          _T_6887_1858 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1859 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h743 == _T_481) begin
          _T_6887_1859 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1860 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h744 == _T_481) begin
          _T_6887_1860 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1861 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h745 == _T_481) begin
          _T_6887_1861 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1862 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h746 == _T_481) begin
          _T_6887_1862 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1863 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h747 == _T_481) begin
          _T_6887_1863 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1864 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h748 == _T_481) begin
          _T_6887_1864 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1865 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h749 == _T_481) begin
          _T_6887_1865 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1866 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74a == _T_481) begin
          _T_6887_1866 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1867 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74b == _T_481) begin
          _T_6887_1867 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1868 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74c == _T_481) begin
          _T_6887_1868 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1869 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74d == _T_481) begin
          _T_6887_1869 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1870 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74e == _T_481) begin
          _T_6887_1870 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1871 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h74f == _T_481) begin
          _T_6887_1871 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1872 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h750 == _T_481) begin
          _T_6887_1872 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1873 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h751 == _T_481) begin
          _T_6887_1873 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1874 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h752 == _T_481) begin
          _T_6887_1874 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1875 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h753 == _T_481) begin
          _T_6887_1875 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1876 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h754 == _T_481) begin
          _T_6887_1876 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1877 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h755 == _T_481) begin
          _T_6887_1877 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1878 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h756 == _T_481) begin
          _T_6887_1878 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1879 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h757 == _T_481) begin
          _T_6887_1879 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1880 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h758 == _T_481) begin
          _T_6887_1880 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1881 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h759 == _T_481) begin
          _T_6887_1881 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1882 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75a == _T_481) begin
          _T_6887_1882 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1883 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75b == _T_481) begin
          _T_6887_1883 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1884 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75c == _T_481) begin
          _T_6887_1884 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1885 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75d == _T_481) begin
          _T_6887_1885 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1886 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75e == _T_481) begin
          _T_6887_1886 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1887 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h75f == _T_481) begin
          _T_6887_1887 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1888 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h760 == _T_481) begin
          _T_6887_1888 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1889 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h761 == _T_481) begin
          _T_6887_1889 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1890 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h762 == _T_481) begin
          _T_6887_1890 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1891 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h763 == _T_481) begin
          _T_6887_1891 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1892 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h764 == _T_481) begin
          _T_6887_1892 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1893 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h765 == _T_481) begin
          _T_6887_1893 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1894 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h766 == _T_481) begin
          _T_6887_1894 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1895 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h767 == _T_481) begin
          _T_6887_1895 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1896 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h768 == _T_481) begin
          _T_6887_1896 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1897 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h769 == _T_481) begin
          _T_6887_1897 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1898 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76a == _T_481) begin
          _T_6887_1898 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1899 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76b == _T_481) begin
          _T_6887_1899 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1900 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76c == _T_481) begin
          _T_6887_1900 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1901 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76d == _T_481) begin
          _T_6887_1901 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1902 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76e == _T_481) begin
          _T_6887_1902 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1903 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h76f == _T_481) begin
          _T_6887_1903 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1904 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h770 == _T_481) begin
          _T_6887_1904 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1905 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h771 == _T_481) begin
          _T_6887_1905 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1906 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h772 == _T_481) begin
          _T_6887_1906 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1907 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h773 == _T_481) begin
          _T_6887_1907 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1908 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h774 == _T_481) begin
          _T_6887_1908 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1909 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h775 == _T_481) begin
          _T_6887_1909 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1910 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h776 == _T_481) begin
          _T_6887_1910 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1911 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h777 == _T_481) begin
          _T_6887_1911 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1912 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h778 == _T_481) begin
          _T_6887_1912 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1913 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h779 == _T_481) begin
          _T_6887_1913 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1914 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77a == _T_481) begin
          _T_6887_1914 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1915 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77b == _T_481) begin
          _T_6887_1915 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1916 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77c == _T_481) begin
          _T_6887_1916 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1917 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77d == _T_481) begin
          _T_6887_1917 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1918 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77e == _T_481) begin
          _T_6887_1918 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1919 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h77f == _T_481) begin
          _T_6887_1919 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1920 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h780 == _T_481) begin
          _T_6887_1920 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1921 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h781 == _T_481) begin
          _T_6887_1921 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1922 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h782 == _T_481) begin
          _T_6887_1922 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1923 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h783 == _T_481) begin
          _T_6887_1923 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1924 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h784 == _T_481) begin
          _T_6887_1924 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1925 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h785 == _T_481) begin
          _T_6887_1925 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1926 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h786 == _T_481) begin
          _T_6887_1926 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1927 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h787 == _T_481) begin
          _T_6887_1927 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1928 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h788 == _T_481) begin
          _T_6887_1928 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1929 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h789 == _T_481) begin
          _T_6887_1929 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1930 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78a == _T_481) begin
          _T_6887_1930 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1931 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78b == _T_481) begin
          _T_6887_1931 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1932 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78c == _T_481) begin
          _T_6887_1932 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1933 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78d == _T_481) begin
          _T_6887_1933 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1934 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78e == _T_481) begin
          _T_6887_1934 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1935 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h78f == _T_481) begin
          _T_6887_1935 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1936 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h790 == _T_481) begin
          _T_6887_1936 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1937 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h791 == _T_481) begin
          _T_6887_1937 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1938 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h792 == _T_481) begin
          _T_6887_1938 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1939 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h793 == _T_481) begin
          _T_6887_1939 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1940 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h794 == _T_481) begin
          _T_6887_1940 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1941 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h795 == _T_481) begin
          _T_6887_1941 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1942 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h796 == _T_481) begin
          _T_6887_1942 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1943 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h797 == _T_481) begin
          _T_6887_1943 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1944 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h798 == _T_481) begin
          _T_6887_1944 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1945 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h799 == _T_481) begin
          _T_6887_1945 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1946 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79a == _T_481) begin
          _T_6887_1946 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1947 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79b == _T_481) begin
          _T_6887_1947 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1948 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79c == _T_481) begin
          _T_6887_1948 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1949 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79d == _T_481) begin
          _T_6887_1949 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1950 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79e == _T_481) begin
          _T_6887_1950 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1951 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h79f == _T_481) begin
          _T_6887_1951 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1952 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a0 == _T_481) begin
          _T_6887_1952 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1953 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a1 == _T_481) begin
          _T_6887_1953 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1954 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a2 == _T_481) begin
          _T_6887_1954 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1955 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a3 == _T_481) begin
          _T_6887_1955 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1956 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a4 == _T_481) begin
          _T_6887_1956 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1957 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a5 == _T_481) begin
          _T_6887_1957 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1958 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a6 == _T_481) begin
          _T_6887_1958 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1959 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a7 == _T_481) begin
          _T_6887_1959 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1960 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a8 == _T_481) begin
          _T_6887_1960 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1961 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7a9 == _T_481) begin
          _T_6887_1961 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1962 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7aa == _T_481) begin
          _T_6887_1962 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1963 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ab == _T_481) begin
          _T_6887_1963 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1964 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ac == _T_481) begin
          _T_6887_1964 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1965 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ad == _T_481) begin
          _T_6887_1965 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1966 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ae == _T_481) begin
          _T_6887_1966 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1967 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7af == _T_481) begin
          _T_6887_1967 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1968 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b0 == _T_481) begin
          _T_6887_1968 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1969 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b1 == _T_481) begin
          _T_6887_1969 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1970 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b2 == _T_481) begin
          _T_6887_1970 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1971 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b3 == _T_481) begin
          _T_6887_1971 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1972 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b4 == _T_481) begin
          _T_6887_1972 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1973 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b5 == _T_481) begin
          _T_6887_1973 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1974 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b6 == _T_481) begin
          _T_6887_1974 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1975 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b7 == _T_481) begin
          _T_6887_1975 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1976 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b8 == _T_481) begin
          _T_6887_1976 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1977 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7b9 == _T_481) begin
          _T_6887_1977 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1978 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ba == _T_481) begin
          _T_6887_1978 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1979 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7bb == _T_481) begin
          _T_6887_1979 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1980 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7bc == _T_481) begin
          _T_6887_1980 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1981 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7bd == _T_481) begin
          _T_6887_1981 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1982 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7be == _T_481) begin
          _T_6887_1982 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1983 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7bf == _T_481) begin
          _T_6887_1983 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1984 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c0 == _T_481) begin
          _T_6887_1984 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1985 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c1 == _T_481) begin
          _T_6887_1985 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1986 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c2 == _T_481) begin
          _T_6887_1986 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1987 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c3 == _T_481) begin
          _T_6887_1987 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1988 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c4 == _T_481) begin
          _T_6887_1988 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1989 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c5 == _T_481) begin
          _T_6887_1989 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1990 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c6 == _T_481) begin
          _T_6887_1990 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1991 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c7 == _T_481) begin
          _T_6887_1991 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1992 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c8 == _T_481) begin
          _T_6887_1992 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1993 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7c9 == _T_481) begin
          _T_6887_1993 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1994 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ca == _T_481) begin
          _T_6887_1994 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1995 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7cb == _T_481) begin
          _T_6887_1995 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1996 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7cc == _T_481) begin
          _T_6887_1996 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1997 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7cd == _T_481) begin
          _T_6887_1997 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1998 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ce == _T_481) begin
          _T_6887_1998 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_1999 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7cf == _T_481) begin
          _T_6887_1999 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2000 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d0 == _T_481) begin
          _T_6887_2000 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2001 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d1 == _T_481) begin
          _T_6887_2001 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2002 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d2 == _T_481) begin
          _T_6887_2002 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2003 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d3 == _T_481) begin
          _T_6887_2003 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2004 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d4 == _T_481) begin
          _T_6887_2004 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2005 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d5 == _T_481) begin
          _T_6887_2005 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2006 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d6 == _T_481) begin
          _T_6887_2006 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2007 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d7 == _T_481) begin
          _T_6887_2007 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2008 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d8 == _T_481) begin
          _T_6887_2008 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2009 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7d9 == _T_481) begin
          _T_6887_2009 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2010 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7da == _T_481) begin
          _T_6887_2010 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2011 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7db == _T_481) begin
          _T_6887_2011 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2012 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7dc == _T_481) begin
          _T_6887_2012 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2013 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7dd == _T_481) begin
          _T_6887_2013 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2014 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7de == _T_481) begin
          _T_6887_2014 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2015 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7df == _T_481) begin
          _T_6887_2015 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2016 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e0 == _T_481) begin
          _T_6887_2016 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2017 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e1 == _T_481) begin
          _T_6887_2017 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2018 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e2 == _T_481) begin
          _T_6887_2018 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2019 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e3 == _T_481) begin
          _T_6887_2019 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2020 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e4 == _T_481) begin
          _T_6887_2020 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2021 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e5 == _T_481) begin
          _T_6887_2021 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2022 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e6 == _T_481) begin
          _T_6887_2022 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2023 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e7 == _T_481) begin
          _T_6887_2023 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2024 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e8 == _T_481) begin
          _T_6887_2024 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2025 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7e9 == _T_481) begin
          _T_6887_2025 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2026 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ea == _T_481) begin
          _T_6887_2026 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2027 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7eb == _T_481) begin
          _T_6887_2027 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2028 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ec == _T_481) begin
          _T_6887_2028 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2029 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ed == _T_481) begin
          _T_6887_2029 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2030 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ee == _T_481) begin
          _T_6887_2030 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2031 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ef == _T_481) begin
          _T_6887_2031 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2032 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f0 == _T_481) begin
          _T_6887_2032 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2033 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f1 == _T_481) begin
          _T_6887_2033 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2034 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f2 == _T_481) begin
          _T_6887_2034 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2035 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f3 == _T_481) begin
          _T_6887_2035 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2036 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f4 == _T_481) begin
          _T_6887_2036 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2037 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f5 == _T_481) begin
          _T_6887_2037 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2038 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f6 == _T_481) begin
          _T_6887_2038 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2039 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f7 == _T_481) begin
          _T_6887_2039 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2040 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f8 == _T_481) begin
          _T_6887_2040 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2041 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7f9 == _T_481) begin
          _T_6887_2041 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2042 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7fa == _T_481) begin
          _T_6887_2042 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2043 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7fb == _T_481) begin
          _T_6887_2043 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2044 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7fc == _T_481) begin
          _T_6887_2044 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2045 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7fd == _T_481) begin
          _T_6887_2045 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2046 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7fe == _T_481) begin
          _T_6887_2046 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_6887_2047 <= 1'h1;
    end else begin
      if (_T_13036) begin
        if (11'h7ff == _T_481) begin
          _T_6887_2047 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_13304_0 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13670) begin
            _T_13304_0 <= _T_13672;
          end else begin
            if (_T_13676) begin
              _T_13304_0 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_1 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13684) begin
            _T_13304_1 <= _T_13672;
          end else begin
            if (_T_13690) begin
              _T_13304_1 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_2 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13698) begin
            _T_13304_2 <= _T_13672;
          end else begin
            if (_T_13704) begin
              _T_13304_2 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_3 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13712) begin
            _T_13304_3 <= _T_13672;
          end else begin
            if (_T_13718) begin
              _T_13304_3 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_4 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13726) begin
            _T_13304_4 <= _T_13672;
          end else begin
            if (_T_13732) begin
              _T_13304_4 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_5 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13740) begin
            _T_13304_5 <= _T_13672;
          end else begin
            if (_T_13746) begin
              _T_13304_5 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_6 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13754) begin
            _T_13304_6 <= _T_13672;
          end else begin
            if (_T_13760) begin
              _T_13304_6 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_7 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13768) begin
            _T_13304_7 <= _T_13672;
          end else begin
            if (_T_13774) begin
              _T_13304_7 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_8 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13782) begin
            _T_13304_8 <= _T_13672;
          end else begin
            if (_T_13788) begin
              _T_13304_8 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_9 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13796) begin
            _T_13304_9 <= _T_13672;
          end else begin
            if (_T_13802) begin
              _T_13304_9 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_10 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13810) begin
            _T_13304_10 <= _T_13672;
          end else begin
            if (_T_13816) begin
              _T_13304_10 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_11 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13824) begin
            _T_13304_11 <= _T_13672;
          end else begin
            if (_T_13830) begin
              _T_13304_11 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_12 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13838) begin
            _T_13304_12 <= _T_13672;
          end else begin
            if (_T_13844) begin
              _T_13304_12 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_13 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13852) begin
            _T_13304_13 <= _T_13672;
          end else begin
            if (_T_13858) begin
              _T_13304_13 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_14 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13866) begin
            _T_13304_14 <= _T_13672;
          end else begin
            if (_T_13872) begin
              _T_13304_14 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13304_15 <= 15'h0;
    end else begin
      if (_T_483) begin
        if (_T_13659) begin
          if (_T_13880) begin
            _T_13304_15 <= _T_13672;
          end else begin
            if (_T_13886) begin
              _T_13304_15 <= _T_13679;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_13893 <= 4'h0;
    end else begin
      if (_T_13896) begin
        if (_T_14097) begin
          _T_13893 <= 4'h0;
        end else begin
          if (_T_13899) begin
            _T_13893 <= _T_14087;
          end
        end
      end else begin
        if (_T_13899) begin
          _T_13893 <= _T_14087;
        end
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else begin
      if (_T_13912) begin
        value_1 <= _T_14153;
      end
    end
    if (_T_14197) begin
      if (3'h7 == value_3) begin
        _T_14075_7 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h7 == _T_14107) begin
            _T_14075_7 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h7 == _T_14096) begin
                if (4'hf == _T_13891) begin
                  _T_14075_7 <= L2_data_array_RW0_rdata_15;
                end else begin
                  if (4'he == _T_13891) begin
                    _T_14075_7 <= L2_data_array_RW0_rdata_14;
                  end else begin
                    if (4'hd == _T_13891) begin
                      _T_14075_7 <= L2_data_array_RW0_rdata_13;
                    end else begin
                      if (4'hc == _T_13891) begin
                        _T_14075_7 <= L2_data_array_RW0_rdata_12;
                      end else begin
                        if (4'hb == _T_13891) begin
                          _T_14075_7 <= L2_data_array_RW0_rdata_11;
                        end else begin
                          if (4'ha == _T_13891) begin
                            _T_14075_7 <= L2_data_array_RW0_rdata_10;
                          end else begin
                            if (4'h9 == _T_13891) begin
                              _T_14075_7 <= L2_data_array_RW0_rdata_9;
                            end else begin
                              if (4'h8 == _T_13891) begin
                                _T_14075_7 <= L2_data_array_RW0_rdata_8;
                              end else begin
                                if (4'h7 == _T_13891) begin
                                  _T_14075_7 <= L2_data_array_RW0_rdata_7;
                                end else begin
                                  if (4'h6 == _T_13891) begin
                                    _T_14075_7 <= L2_data_array_RW0_rdata_6;
                                  end else begin
                                    if (4'h5 == _T_13891) begin
                                      _T_14075_7 <= L2_data_array_RW0_rdata_5;
                                    end else begin
                                      if (4'h4 == _T_13891) begin
                                        _T_14075_7 <= L2_data_array_RW0_rdata_4;
                                      end else begin
                                        if (4'h3 == _T_13891) begin
                                          _T_14075_7 <= L2_data_array_RW0_rdata_3;
                                        end else begin
                                          if (4'h2 == _T_13891) begin
                                            _T_14075_7 <= L2_data_array_RW0_rdata_2;
                                          end else begin
                                            if (4'h1 == _T_13891) begin
                                              _T_14075_7 <= L2_data_array_RW0_rdata_1;
                                            end else begin
                                              _T_14075_7 <= _GEN_6883;
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h7 == _T_14096) begin
              if (4'hf == _T_13891) begin
                _T_14075_7 <= L2_data_array_RW0_rdata_15;
              end else begin
                if (4'he == _T_13891) begin
                  _T_14075_7 <= L2_data_array_RW0_rdata_14;
                end else begin
                  if (4'hd == _T_13891) begin
                    _T_14075_7 <= L2_data_array_RW0_rdata_13;
                  end else begin
                    if (4'hc == _T_13891) begin
                      _T_14075_7 <= L2_data_array_RW0_rdata_12;
                    end else begin
                      if (4'hb == _T_13891) begin
                        _T_14075_7 <= L2_data_array_RW0_rdata_11;
                      end else begin
                        if (4'ha == _T_13891) begin
                          _T_14075_7 <= L2_data_array_RW0_rdata_10;
                        end else begin
                          if (4'h9 == _T_13891) begin
                            _T_14075_7 <= L2_data_array_RW0_rdata_9;
                          end else begin
                            if (4'h8 == _T_13891) begin
                              _T_14075_7 <= L2_data_array_RW0_rdata_8;
                            end else begin
                              if (4'h7 == _T_13891) begin
                                _T_14075_7 <= L2_data_array_RW0_rdata_7;
                              end else begin
                                if (4'h6 == _T_13891) begin
                                  _T_14075_7 <= L2_data_array_RW0_rdata_6;
                                end else begin
                                  if (4'h5 == _T_13891) begin
                                    _T_14075_7 <= L2_data_array_RW0_rdata_5;
                                  end else begin
                                    if (4'h4 == _T_13891) begin
                                      _T_14075_7 <= L2_data_array_RW0_rdata_4;
                                    end else begin
                                      if (4'h3 == _T_13891) begin
                                        _T_14075_7 <= L2_data_array_RW0_rdata_3;
                                      end else begin
                                        if (4'h2 == _T_13891) begin
                                          _T_14075_7 <= L2_data_array_RW0_rdata_2;
                                        end else begin
                                          if (4'h1 == _T_13891) begin
                                            _T_14075_7 <= L2_data_array_RW0_rdata_1;
                                          end else begin
                                            _T_14075_7 <= _GEN_6883;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h7 == _T_14107) begin
          _T_14075_7 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h7 == _T_14096) begin
              if (4'hf == _T_13891) begin
                _T_14075_7 <= L2_data_array_RW0_rdata_15;
              end else begin
                if (4'he == _T_13891) begin
                  _T_14075_7 <= L2_data_array_RW0_rdata_14;
                end else begin
                  if (4'hd == _T_13891) begin
                    _T_14075_7 <= L2_data_array_RW0_rdata_13;
                  end else begin
                    if (4'hc == _T_13891) begin
                      _T_14075_7 <= L2_data_array_RW0_rdata_12;
                    end else begin
                      if (4'hb == _T_13891) begin
                        _T_14075_7 <= L2_data_array_RW0_rdata_11;
                      end else begin
                        if (4'ha == _T_13891) begin
                          _T_14075_7 <= L2_data_array_RW0_rdata_10;
                        end else begin
                          if (4'h9 == _T_13891) begin
                            _T_14075_7 <= L2_data_array_RW0_rdata_9;
                          end else begin
                            if (4'h8 == _T_13891) begin
                              _T_14075_7 <= L2_data_array_RW0_rdata_8;
                            end else begin
                              if (4'h7 == _T_13891) begin
                                _T_14075_7 <= L2_data_array_RW0_rdata_7;
                              end else begin
                                if (4'h6 == _T_13891) begin
                                  _T_14075_7 <= L2_data_array_RW0_rdata_6;
                                end else begin
                                  if (4'h5 == _T_13891) begin
                                    _T_14075_7 <= L2_data_array_RW0_rdata_5;
                                  end else begin
                                    if (4'h4 == _T_13891) begin
                                      _T_14075_7 <= L2_data_array_RW0_rdata_4;
                                    end else begin
                                      if (4'h3 == _T_13891) begin
                                        _T_14075_7 <= L2_data_array_RW0_rdata_3;
                                      end else begin
                                        if (4'h2 == _T_13891) begin
                                          _T_14075_7 <= L2_data_array_RW0_rdata_2;
                                        end else begin
                                          if (4'h1 == _T_13891) begin
                                            _T_14075_7 <= L2_data_array_RW0_rdata_1;
                                          end else begin
                                            _T_14075_7 <= _GEN_6883;
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h7 == _T_14096) begin
            if (4'hf == _T_13891) begin
              _T_14075_7 <= L2_data_array_RW0_rdata_15;
            end else begin
              if (4'he == _T_13891) begin
                _T_14075_7 <= L2_data_array_RW0_rdata_14;
              end else begin
                if (4'hd == _T_13891) begin
                  _T_14075_7 <= L2_data_array_RW0_rdata_13;
                end else begin
                  if (4'hc == _T_13891) begin
                    _T_14075_7 <= L2_data_array_RW0_rdata_12;
                  end else begin
                    if (4'hb == _T_13891) begin
                      _T_14075_7 <= L2_data_array_RW0_rdata_11;
                    end else begin
                      if (4'ha == _T_13891) begin
                        _T_14075_7 <= L2_data_array_RW0_rdata_10;
                      end else begin
                        if (4'h9 == _T_13891) begin
                          _T_14075_7 <= L2_data_array_RW0_rdata_9;
                        end else begin
                          if (4'h8 == _T_13891) begin
                            _T_14075_7 <= L2_data_array_RW0_rdata_8;
                          end else begin
                            if (4'h7 == _T_13891) begin
                              _T_14075_7 <= L2_data_array_RW0_rdata_7;
                            end else begin
                              if (4'h6 == _T_13891) begin
                                _T_14075_7 <= L2_data_array_RW0_rdata_6;
                              end else begin
                                if (4'h5 == _T_13891) begin
                                  _T_14075_7 <= L2_data_array_RW0_rdata_5;
                                end else begin
                                  if (4'h4 == _T_13891) begin
                                    _T_14075_7 <= L2_data_array_RW0_rdata_4;
                                  end else begin
                                    if (4'h3 == _T_13891) begin
                                      _T_14075_7 <= L2_data_array_RW0_rdata_3;
                                    end else begin
                                      if (4'h2 == _T_13891) begin
                                        _T_14075_7 <= L2_data_array_RW0_rdata_2;
                                      end else begin
                                        if (4'h1 == _T_13891) begin
                                          _T_14075_7 <= L2_data_array_RW0_rdata_1;
                                        end else begin
                                          _T_14075_7 <= _GEN_6883;
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h6 == value_3) begin
        _T_14075_6 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h6 == _T_14107) begin
            _T_14075_6 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h6 == _T_14096) begin
                _T_14075_6 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h6 == _T_14096) begin
              _T_14075_6 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h6 == _T_14107) begin
          _T_14075_6 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h6 == _T_14096) begin
              _T_14075_6 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h6 == _T_14096) begin
            _T_14075_6 <= _GEN_6898;
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h5 == value_3) begin
        _T_14075_5 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h5 == _T_14107) begin
            _T_14075_5 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h5 == _T_14096) begin
                _T_14075_5 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h5 == _T_14096) begin
              _T_14075_5 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h5 == _T_14107) begin
          _T_14075_5 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h5 == _T_14096) begin
              _T_14075_5 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h5 == _T_14096) begin
            _T_14075_5 <= _GEN_6898;
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h4 == value_3) begin
        _T_14075_4 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h4 == _T_14107) begin
            _T_14075_4 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h4 == _T_14096) begin
                _T_14075_4 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h4 == _T_14096) begin
              _T_14075_4 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h4 == _T_14107) begin
          _T_14075_4 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h4 == _T_14096) begin
              _T_14075_4 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h4 == _T_14096) begin
            _T_14075_4 <= _GEN_6898;
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h3 == value_3) begin
        _T_14075_3 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h3 == _T_14107) begin
            _T_14075_3 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h3 == _T_14096) begin
                _T_14075_3 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h3 == _T_14096) begin
              _T_14075_3 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h3 == _T_14107) begin
          _T_14075_3 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h3 == _T_14096) begin
              _T_14075_3 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h3 == _T_14096) begin
            _T_14075_3 <= _GEN_6898;
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h2 == value_3) begin
        _T_14075_2 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h2 == _T_14107) begin
            _T_14075_2 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h2 == _T_14096) begin
                _T_14075_2 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h2 == _T_14096) begin
              _T_14075_2 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h2 == _T_14107) begin
          _T_14075_2 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h2 == _T_14096) begin
              _T_14075_2 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h2 == _T_14096) begin
            _T_14075_2 <= _GEN_6898;
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h1 == value_3) begin
        _T_14075_1 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h1 == _T_14107) begin
            _T_14075_1 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h1 == _T_14096) begin
                _T_14075_1 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h1 == _T_14096) begin
              _T_14075_1 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h1 == _T_14107) begin
          _T_14075_1 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h1 == _T_14096) begin
              _T_14075_1 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h1 == _T_14096) begin
            _T_14075_1 <= _GEN_6898;
          end
        end
      end
    end
    if (_T_14197) begin
      if (3'h0 == value_3) begin
        _T_14075_0 <= auto_out_d_bits_data;
      end else begin
        if (_T_14102) begin
          if (3'h0 == _T_14107) begin
            _T_14075_0 <= _T_14148;
          end else begin
            if (_T_13896) begin
              if (3'h0 == _T_14096) begin
                _T_14075_0 <= _GEN_6898;
              end
            end
          end
        end else begin
          if (_T_13896) begin
            if (3'h0 == _T_14096) begin
              _T_14075_0 <= _GEN_6898;
            end
          end
        end
      end
    end else begin
      if (_T_14102) begin
        if (3'h0 == _T_14107) begin
          _T_14075_0 <= _T_14148;
        end else begin
          if (_T_13896) begin
            if (3'h0 == _T_14096) begin
              _T_14075_0 <= _GEN_6898;
            end
          end
        end
      end else begin
        if (_T_13896) begin
          if (3'h0 == _T_14096) begin
            _T_14075_0 <= _GEN_6898;
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else begin
      if (_T_14172) begin
        value_2 <= _T_14176;
      end
    end
    if (reset) begin
      value_3 <= 3'h0;
    end else begin
      if (_T_14190) begin
        value_3 <= _T_14194;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (1'h0) begin
          $fwrite(32'h80000002,"Assertion failed: Inner tilelink Unexpected handshake\n    at TLSimpleL2.scala:239 assert(N, \"Inner tilelink Unexpected handshake\")\n"); // @[TLSimpleL2.scala 239:17:freechips.rocketchip.system.DefaultConfig.fir@221116.14]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (1'h0) begin
          $fatal; // @[TLSimpleL2.scala 239:17:freechips.rocketchip.system.DefaultConfig.fir@221117.14]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7036 & _T_261) begin
          $fwrite(32'h80000002,"Assertion failed: state error\n    at TLSimpleL2.scala:260 assert(N, \"state error\")\n"); // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221170.12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7036 & _T_261) begin
          $fatal; // @[TLSimpleL2.scala 260:17:freechips.rocketchip.system.DefaultConfig.fir@221171.12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_482 & _T_13388) begin
          $fwrite(32'h80000002,"Assertion failed: cross cache line bursts detected\n    at TLSimpleL2.scala:395 assert(inner_end_beat < innerDataBeats.U, \"cross cache line bursts detected\")\n"); // @[TLSimpleL2.scala 395:15:freechips.rocketchip.system.DefaultConfig.fir@223722.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_482 & _T_13388) begin
          $fatal; // @[TLSimpleL2.scala 395:15:freechips.rocketchip.system.DefaultConfig.fir@223723.8]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7044 & _T_261) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected condition in s_tag_read\n    at TLSimpleL2.scala:403 assert(N, \"Unexpected condition in s_tag_read\")\n"); // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223741.12]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7044 & _T_261) begin
          $fatal; // @[TLSimpleL2.scala 403:17:freechips.rocketchip.system.DefaultConfig.fir@223742.12]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7049 & _T_13663) begin
          $fwrite(32'h80000002,"Assertion failed: update must = repl way when decrease a dsid's occupacy\n    at TLSimpleL2.scala:462 assert(update_way === repl_way, \"update must = repl way when decrease a dsid's occupacy\")\n"); // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224190.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7049 & _T_13663) begin
          $fatal; // @[TLSimpleL2.scala 462:17:freechips.rocketchip.system.DefaultConfig.fir@224191.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7057 & _T_261) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected condition in s_data_read\n    at TLSimpleL2.scala:532 assert(N, \"Unexpected condition in s_data_read\")\n"); // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224702.16]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7057 & _T_261) begin
          $fatal; // @[TLSimpleL2.scala 532:19:freechips.rocketchip.system.DefaultConfig.fir@224703.16]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_7066 & _T_261) begin
          $fwrite(32'h80000002,"Assertion failed: Unexpected condition in s_wait_ram_bresp\n    at TLSimpleL2.scala:602 assert(N, \"Unexpected condition in s_wait_ram_bresp\")\n"); // @[TLSimpleL2.scala 602:17:freechips.rocketchip.system.DefaultConfig.fir@224821.10]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_7066 & _T_261) begin
          $fatal; // @[TLSimpleL2.scala 602:17:freechips.rocketchip.system.DefaultConfig.fir@224822.10]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
